// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:07 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rBOQuf5Ykl+Eluc/U+ii0HgPPPADt0vmaZg4TWpc2W4cHWkQ6u+rwPXfp309uCCy
IGZBjjCWeWE7f4R9fsvsylS4uLA9a4BrCBq48c2nW0gd+52h2AfdTYcM5G2Kj8SO
Y92lm07cDiTl0+JKqYngYr78sECDW274j6ipZe3RBcM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
XVg+a1SxKGSPJQFuibB1dmGdzpLvLSdSHWLXmE4PMVlZu5ed1t6JUF9yoNhsJolj
JaYlVUMjVw/aNRDB7fUzAYNWdYoUwblujDjBxwado2KjEiIvqd3mU3kYSUCjgiIp
NOr/bdToFPmvaEbHlGxhVJ4eK1L8fY0lL1HkuYUqTDl2RPDjBlTWHtx7YT/hhWhZ
snpVd+cAQDgxQDyS6dC7+1dFW18izSiffwiFljMlz3SftxMYsrgtg0sQ/IIkNeDQ
aWlCuwXYtR0uNR9Tg3qj7Fr+nUpZXtG4lksksK0Q21aobwUhK5hV7rzSHSbN1YzJ
QKC9QmutANfIkpfc8Q4v1TmqTwao2YaKaC3ql8mYWbbguzAcXrg7R9wtvgxihZdR
mrOYsWq/4vK7aHe4PFa4taGPNuhufOh45KF6bJwDd5n+gc+hO5PDlScCqNOYFYy/
aldWOFeMILyNdPuHJ+NDz70EYD3+4ZCiaMfHjS2c//+fjJnCxUTmdr+KsPaMoJwS
FF7dfKWqZSMjAyJn+ScHpDQs4mBDAeIN0y2LmJDkhmkdhlFFk04LNP7ZNQDUksm4
qRJh3rrP70UJk5VdcpRygFCW1kgramWuxo1AL5cxlWbyPtjOvcSJpdaRWFb1O+Dc
CPkwRq1GwNgMeXkUz1aCxKQ4/8ivGERCZ0czqZW+egTNa7gZQV6k8ZLhFo6Tc87+
DH6G+C6VGKhk9GoT13FmeWj1pcfLuwvJJUfZ2c9seh9nUH0UC6glrOVvbMRgi1I/
JxL5tWBFtqIH22fusj9jGT7BOZdaoSDh1DXgLP1moArR9n4pGNwKXyp3r5/a1KZw
WUREBJp/lT73rgwX/+p0U6o+yqkp/gi37b0g9X9bA1yMV1lrBdVSS/7n3eq86muB
016ipwde0+W4mJ8Osc1jI96b+68ripkkl4OxikNYe8n2pU67P1hl7bLDc6IC8JE9
u0+t1rlEF5mQyyZEUz5d0fmJTEtBUGwnt35fpbh0bXf4jbDyX08NULIhbi95EcTD
QZ9YF4oiSsNceac1RJZuJezJaF7zSJS0QMa3gKLoZcYvr/YvbX8b7FoCf4hNualm
IjD03xb/uloWNyBpHrNKNecrexsuYDVvWn7bTi/PrqeiJlaPeIWO62mM9nL9jswX
8AM4n4uzXst2x+gtL9r2fmnwX/on0Uc7LgsB2fabWPhT6hxFt1DeIQ7oTz5XxWx1
AlPCBVA7lmA5YabAVvy44HiF/9tLewGS+id3qh2wUPCOsy5SAVsoxmPBxPVscLjm
2cxpEpp+hPgbUlLnV5pJa0f82O+khtw9UUKqusT+kBlXpu57BPhLC5biu/793XdB
wDSF9KCj2t6G0J08ozSIwW/Ev8nX01MvN5DTHVklgub3Je1F4Q/2QSUI0vWFGr61
5cUi1BVf08hKZXYGYbHTTO0JizjFZ/ay6UpQMiFQVOGFa/rEoQakAIHGZlTGWW6Q
ofMAQSw2sdnUPwIEljr2mV/UsAoUJHvJw+Grgg6r7c7DTl7KomdZ32XbUBujXYSW
/a2ReHcjhhWVMQTCqROaZJjWreeAULJ0xLRfDuy24mL2Qj253qH97tLUVM0KlGro
XKSty6kl43q9g4LdbQrtAoeKyHy63Ml6vciDuFxFKv+Cm2+H4mmnVWzKCr09Skls
DSb9DXQGojSC09afhwWpnmaelS8GzUTsvXprtFQWgFMuDTUWZ4X6ypurhW2XdVpO
LE6ZC7dekHXvAldTpHbkY1W3MNUvcNBNb3YOGecQS2UxVGPqJ7tiBwJDNSI7t2al
FEqJBwLB0BwJCDVkWOdqRvEZH8Uo8igFFiJgGcfmq7/3JgvPSzEePU8JfVYY1ZsK
e5CDyYqRIPv/UOuQmWbE03lA1MC9Pb5pVlPMDolPtidZgiYAPVDEgQmK/w8v3d7P
D5gq1tOtwX3vkuZBAsegPzbxIZl7QIfOs82QIif3YXo+Zwb5RPB8PBua6n4Fn9RQ
G/DdQjcGPlhteW3IpKZipAbqsUy1opY7De8/BK9nmHl5hn/kbWQq4gpIoPJzKALX
v+s+1JMOpANZyQDRK+1/wsH4LVh8hBL3Jj3hA0X505g4dU4riTHefNakVBHUMe3l
iMgbgQ/dpkOdwWchcbkFNfXg6pfYzLkVpYTHmVy4OyY7CnwwM3DVIFEr1j9aGXfR
pvQbw6UubIwnVRCBtGWOkTHnY7QD1eGxSKaKYYzDX9JjuuWyZQC1pv7nAfqX0EKb
jvHeklI5rWSz7jhnACIJs1EmOxaifpdROFmZiTALUmZUMz7dEbwMI6iATOhYL8oe
Xs4tZuZDYx75sO4cM/hBYYhbYkiD5jCcc3cDNzn8OX80eyA4hhPXLGRL218Ov8jp
06bpTQtWzz08bfGr0KXhQqdxCPiYLlsuCp42WOG3QkVsrALQbRAuY/iTDvJ9xU8Z
okMOOFpxzgvMweibd7zUyzZRGIOFsmFV8kiFnD3ZewApzPsX3GGHnRPOEfhEfnqj
4ZDl+BBfV5E5V5t01L+yUlYHVqTbtUfv4Vqy6XFub/ffUOfxwInls9os+V5feksA
kX8lJKU3AYWKBM7xr+4gvSodKfxDRy/vJtk4JlVs7yPTKtbpQqP8/PgCgAXpXH6K
229uM5p4BVyxLFMPvIasGDVQLLBQ2NGCeq3G3h2wSRPlBXveWiIddaBb4k5oZHJ1
7rwCE5YHxBOVGfNuIKw7ZJQnz7/Fy72k+flVb+eRcAPDaiAPI3k99eoLKN3VOaR6
ZuTtdN1WRiT3NAatVYmK+CJEcHi1P9XevsxhLF7B5F6zYwNXsaLK2l4bw5tBYA1a
MBfloDCzal7Yu4qOhikWFGRmLt2VMj+Ove9yAZX6i+l/uaDsR5vjb9Lkp/oQUZw3
88ZZ9vu4tBecj577QhpoL74YT/bc58dvPA0hS/LoOiDGs4Jo+Hh1UQoq7uUz1v4H
sjL+2gaGLrmtLWRLbALu0KoCS7kUId+17io4altaP2kVdCZqKG3esWStHwgrABx5
UiTKWA+K0jdwZOYbbv0ZEFlpAccY9TqezKuFdIwSEP+koCtjKZiyH89RIlZ1OmBt
x4bSFaMFzbe2Ul1tIc+WDesPJE/m4ZOM6xiXAFyDUYTHrmKqtu3tUaCFudWrZmit
R0FvFABf6PGsp0P2Iu5F7p9cXVLDkqrJSbiOBQeshw24SzRUvRFq1QUTPlr1BgLT
ONouVPEbdWikmdnYRNLO3Aydb7uXr1UjGA7fhrQXFhZqEiGp0XoDVWbhVmQZQTSA
EoA77vSZGibgNu5Z4Wpm2zJV13uQI97IL7swsnRPrssLUlCoZl6hZWUL1ZIryFet
ZleLC3xK1OT77AgtRXxgS1f+VmtwG5ZTjrcVfP5PvMdOXvIuHg6VezVPiwtNc0Wf
WNxPoPtI3C5IPg7UJ0eAW+zYSDwETF3sM0/tAumlQUHO5gNFxOgv1inT1oJ+8J3W
Z4JDVwHS9k9X57SVoYn8GVN3zbdZADCm3Cx8OFgIO90yqGXVb1w5SZjUI64sVpSX
16kohnsHbhZIZJGuXkQeUt6x0Q6JsjFDhGWPIRks/hAOVJCZvUKghhUwiGjOHJLR
9UzdUyEL81IENQClwTcz42aYH8Ihf9s2XeoU1y97vZHK8MmtPTlGRwvYOkCRflEK
CVy/nk/vyE5uZ4gJ4gcM+4l/UzlYlXr1TuhM5GxbXxFSHpi7yOjFvriLdOwOu4L7
X5aRCOKgMcBcQUIuBdalOvFiofT1E4mq8qTj4Fd119eJ0bodiI+Apw8JZGMHz2Cl
q8475mHfwZX+OghXB7UsavB9lPOKvz2gVBQbf9sPyWXcs7lhzaBIOWphRhCbOQ6D
K1NKLLtmZrBY/Sf+nZEmE8bh7j5BSzrq7QpIVApOJZPgQBrdnX25sKmBUXW0maW8
RVLQJUNYNSTfsEeEWXIKjG/JCTHPYHt6Y/tySfObt6fqUDBU/JzkbSdOjcFF6WlK
HM0VCsB8GVCd3KjbzJipOw6oVhu3KMFMqK/IPWRDJce2K5K07gEjn6U8LQ6S5M8c
8/PNXXaUmij7JcLUoP/s6OPjOK9zwXoALM5Ot7EZw1FSfkMQ56U67shuXccCg0iy
v6zT1MKJqosj8WWfjglIdSU/w4V5tt+7ZHMXY8FufmhG2LkfHvpYJkgMvtuGpf2P
DIezJmT8GsdXRaWOVM4nyPIf6GVkT9owu4E21ESXWQ34w24r5XzbNy3RSgjRxXK0
9l6JosVulNfkVHm4pFzt3YY+9QiYmjbysJjSjjlZmpaR95y7iteALpkpjjMOeocZ
OwiC8bzQi4/uzzd4xr8puflaTEiaYUX4/Zw5Wq3OdWQlG0/0ddkz4Ow/hNzqbrU0
5RX18a6nZcHeSiRuCp8FH9ZSwuX+3q1qZsa0HJEXVmegGNqqee9kUqk4R68iIyYG
Sq+Jam3cCSHTg114DLHEEU/+5M3eT1aLEhdSPqKNcUJsVUToE/MGq0JQaxpg3u3b
TFFZVBg6YC6OeZnS8EeGXf+97D8C0nsis0sXlvfamY8pmqu4WjRqi36/Mj3Q2FfG
GyoGtNI11xUCbea05v5FjrR90VnIY2CW7bKiUoqbRIgvhFs6ITvM/FIKOoOJfNKi
hswsf4ZK46oe6n8I4NZX/IyYb4abPRVRXa6q5OkL8FhVhl6jL2fKhbIAc02HOWk7
URR6+IB9ZAJtYlyjGfMe03SSo9QeVnhJYDKbjWwdGwaCrbHDPVPORGbb7uI3UsYX
fguXEgpIBr+1avqrjZ6mx0nGrMl6Em7RHbjzA/iqm7lKYkmtQM3sZ96SvOKKRnpu
4MeJA66C535HRbC4nvrqH4N8sWjFHqrfs0iMlf7ANnLzsFuC06D4jTOoxTaeRPxY
7qMigIHKW5iNZ+oCjfpsCHPaRXCn4AuZyAA6A4eLW74fwhYDuF+wF3NllGfsoA/w
lxFAKzDwf/HMc3Zg0sUbUod25fFnL0DPGPcK7C4b0EY6VWg06SGZNjTr9Hbd/XdY
2ax/sKRHF2tvIt7uD76tTjm1IPq4OMpZuJJ9oGSN+5JgcM+TE9y3ZoC9GztcVqGT
lqIDJ5RX8lZr/CeNOVwQieZpDM/HOLVEXUnno7WVuemHTFFg00EGUtTsiVoAr6Vd
nAL8sZ8ctO0OfQkH/GeTUPSaBVs3ZzW7b3XHoR7HpA5pi78KuKkWuhx5GHG7dx3M
uSZYCnulN+nDhYngpgE6NgEdy5hmTYWx9gajZsnZx7mTP4RXhTJp2wl28EHgme03
JSd1SpB6QF7ov2RgVLEI/JtgToO4mJt2Jzh9LxEctkbB9DH83mDMuXGklnGZB4V0
1Qaya6sXRjJ2p2efysG00vXjlVhGYhXLHGYJgQOnbnDWEuqWzgr7vBdlVJVy1ypk
heU9V1OiyFvdsSY1IcLXje8TQF8kF7259mzXipZnCUNjvLSI8Paca7LfBlN9BoAv
lOA+U1uB0e+q6QVrNUVlbrwzJvAcgq7Lo5qDLvaMTQkk7M7tOhCapf+0+lpdIUbi
L+2jqSII9zvWHb7BzXqCA4krA+rIW4z6+nshv5Y2mbauUgEXt6xDYFuuQlAwHJnm
NXLnxV7yhSenBUoAzn5vr2H2rbXjFmiroMLengxiluodGw+qCpQZiRKGZ80UmaIi
IuRXoMzR2f/8EzVUs0d/VisO2HX+GOCfwbTev9nGH0RaP071QSyt9N6vCd8Theg5
Q1F5jT7VVf7+yOekY/pL9LucmNKHYljKDa5pQ/0+0MJIBCksXWogCGAGCYN8MXkk
GFJZlX6LEqfJ1RqU0wDMDFBmal+XV5TJ4aFusrLFnz6tW6MhhGd9OHFH79Ni5kbv
c6qJswW56NPaltMnreeHuIJfA0RvLW31sW4pXLvsPSg+fsRqg8ghcD/geFMvlZ0g
YjRhys0gcnCMYDoBiUF6+wBH+iZ1bvlaVlmkWZmMidya0IvvGHtE/iIGcN1yToiI
yo1Q6Yn2q+zlyDVNfyaiDPKSnrI3qSiR6ghPfwn2/IxzlBBx83fRHQ3MZSliGRqO
wmkRkchuTVsP9jyqB5hW/R820/uPxRxbeHgX1nqJuJkAHbacCSiNqcUapPNJMfz7
+wPusP+TApNF08v09mRWbWs+XXaqMyBju4rTjBtBjnXrVh26W+A8t8rGVEjhCo8+
Ig6Gz+/XTBu9VK8oNG3WTpvaIrukZmUsYoFFAVytqN02Ln0j1RoFzs1BezYoxyvw
jToV5FaZe/QATK0RVIh2wDpClhVL7xaF9nWBMEoZREqb4s0o1xZ/q15ylPwR5qfk
LjtRgA1YEMjK0zDjB9Ppeqd8eIl4Ftrt9V2p0f4bpeGgX+5wrKtP5OIIIP6BcvOR
KJYI+Zyco62K6NHsGQItuQfTNy59sq954L5AOKcx4Aj6HWiw9Twa/R4uBhj6eAZE
eHnzg0ypUAmZAApeCipuOVjv6KO7ZW3Cdq+fXsKrcc5R8io1oeDmTu8wgOeYQgSE
l5jCvPCrpjFhtVxgNdRcAzQrffEC9YHDNu3InCpUJJt8lr6MYH+Kcphr+27K6f77
WHc8vhQF4WA7tq4+T/YiAEdiy7AZgpNqLp0iAWRQXNfx4lqOwDMxq4Hz9eldjipw
fu3jFiZQmpitM+lGmbuxNKu/RtJ2z2kFhT/fwbLqZv5z1HjEWWCp8eqyHmhozFFC
8m3p1QVEDOmb0RYVz5B8myKv7Jo7BDQXAWISdwtI38bRMjyHZheMdIwoMQJ4TaiP
SRL9yHfUlV45/Sfeg46Wu8vhBGbKNUXFFxe2o07uDEl+naYMZobpJD329a8M416t
6kjNvT3b2VIePzl5KVQBs3+fe7HwbkTn24REhYXC9UdpGtsqhalWmOon4SXdgDMs
bJJs3hR3JlRqKEw/DEOoK06BFakkP1HcVJB9k/ECa92MNBbSuoqMvjfn7HsqoTmj
SOtJqLNY05PCOHulYduqUEvV5TYhMIb4Vg4KtzrrvJSjy9A4rHJJzo6JoKc1e9/B
uWNqW4JXwmHalWPH2fqOn1RnI/cGAM4pAHeBAbQ5sbc3EvhVJdeld23yytZHeQFL
nWfN/xcV9qUn8whDWKbhjaqlVJvdI3pa+xDQljNSTB1RhVGniKUUUjMpuxu7FS+Y
dbBdlpqXM2Rt1kHQFYE0CGelQerjT9643KKzXqu9Fa7DHS1J25q0DRsoaibg3LEo
Qwh55AvO0O8GZ7E0FkgmFe/nJGcgFE1wzjz4MrQriyyzgHbmT4WKzUOF+azREZCp
QJwIB3qa9ZuCO7B3lxibFEHlAbSO1kb+VwYLGeHJtbUUKv4650XZo3g9dgo07M3G
YeqHQ4wTUVsZAYC/NfLYYVp3y8wh4vRpT0ZvvKHWRHfyKMd3hCYPDZs5sNXbYOjJ
dLhlpwYd/KUyCINrQfmH8LVb8T9Xh+Q8mWcZ7AChlHGb1eGtKwttSF+MSSwC2wil
zOS9N4079BmG2fP8Q5p/qQmWnReXqbmuXjFgG1cKrrrtnkO8Y0e9rSEMtFQwbH7T
i+PE0TjUxWb3UjT4efxwQksY/eziq2EdB1sust4G4sz4TDFw+ewbpFA4TlJpr1yA
hHVqEpEs3xwa47SlR+Cl0atj20Ir03uknzskIDUvxBuQbsglse7K+W9FiqtCIE9S
veiq2N46FuqGLzYf4GD+Ygopm7qeJCLD6XuU64RqGMF8Uxc+wI2Mkzovg/mzTGbo
xlJV+yKfTYB8X3kIQkWvr0xn3Vu9qXWsqlhwQNczRezIzubBu/eS/7a6MFk+gew2
j7n/WL0LTawv9TuvfJ7XiqE24kqbqnmaEH6TfP91BK87lY6zaKyOl1Mm3ycpU2ov
7CcWZ597AZL/R19tJfXcl2couxPWiIhQb4vMUsIJRyR4+qvulyOoYdwk0OW++uqr
Et8IdJeJn+d8m9JeBxzBZwa0qKi+V6iIgi07BZ3VaOytWcPMBr+JQ+BjK7daaZDv
iDxmHNr2ww4QHoH0CWbHm3KbAj2DyN6GuqcppJcJobFbKAywcpnHzzRK9+/o4Vxd
rrEvqbRH/wnvaKWEA4ZKye6ndxCK6RplvKHfD3uCNbWuIFV0VaI6O3h1QXWCh3DY
+JNBpOvzt/djnc5KK2gkqQJffzxggzIX4w6Ta1VTg42Y7BFIBy+/yeQrS83ZUN0R
Nec2CvndOrNX6ixtD5B89QdzWTNAgKXq20g74xKvA/vTXp1P1KbZTIxfwfURYW3l
y9O+yKkDnSz0Ml17v7E4HZPw8g+j2G4TvNxghf6sZPpd+8fnOPsQHI8T18TYFazA
Vvl6Ei79PibYqE+ET5luRyMUmmxc8dvI4ggfLGWewH/07y7RJpFJ2fFNIGKfX3KQ
kMLVVeCqzNrvG0Wtyc1Eky2u7EhzPhKT5Y0WgzLtMc+q3SfnXb72wkfnwzS9hlUk
wXLxFaLFYYZosBXIJjCkNwXPzZsUdX+bGx7deUzTg9Y4pH0ZIl6ShlqjQTny0gBr
M4Fk5XmVv533sLAtWWwB3VZu8VTkRVAGF7Kml78JapjD+gqhY02+95zySESK5Zwz
M5XdWILnK3HVsxzpMfNSdA==
`pragma protect end_protected
