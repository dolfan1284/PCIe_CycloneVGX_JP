// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:05 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U9/DWMpTN4ws054oYrwoO/lkOcgZUKJTdIBsy5GFTA5NpHI2G0PZNuFlQWGkt842
xmqvZZiX7QRf93+9jNhqI6nGNwnbCg6ZpNeJ5DU54SRzWulVWVYvWm/0QbwAoS8n
64JVPpBiWm/6OwzoyvHm4RPZfgQ97MB9sV6bQO2rD14=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
n2tHr+GPyfUbiuy023wbiiJLAUXCVw0axqCZemWnCvIWLYxpqGLoFnApn4LQHk6A
scgppdrJffsxlwOSfQqBDdXBCVLSDCC0834Tw2kcnoFFOdkkNEqM/W0pmU9hTb+a
7zUg5BkOO6HvNdQG0LMDjpnA3XcYxztuKArh21bKJojVG8gb3gy0b2lvtxiUQjsw
ouGjCshAvFhKxkJpvtR8bh+IAln6WdjOacv58YHedabUzQ0AGddYGT47QYLJQo+o
N1IidM3iJDVelVg40ZgCxpfXpbftsyId3FnOG+k87ntMdZbJ6fJQSdMHR+7e+gxD
bEKSpfHJDrUmdYT+VMEVHaMvFBKCHEojXb8g5xQ7VZcE1cvjOoJHX0cJdJ45HRsC
5SHBIFyifJBsZsHgV6t2pNBlM/kay1bkUy3Hjf18hWKjpE/Pc51CqxngjknPkrAT
XFPfUAY+K2lnFqVU9QxRbMPhZgfgi7z9S7l72xRUyDTZd5o2fhQi9nroOlKpyq2E
XAEnHR2ahQDmNEDAZN22XrHfnKNoTR85Gel6Wmr1FYCMBp1TDfj901HZ8ouQ7TDF
bnS+DSJkE6suWvAAZCTFtum/sHLx8kIbxjVA7dzjTRbxa934fTLZBtD11wvjZVRn
gmoqzseNJBcJhHaD/16NzAb7jWctDLOJyCA3iVbkkZz+D4tV0Xc/QuEbHTEQlpvy
Qzu6u6DFfjAv+m5lNOhlNRiz4LElodPA3/7LCNnoezEvH5LrQNyxIf43sPssUak2
fJkdCCtnh9VaAwk2hiPomf9zq0SueOoz2TqiYHOfyrbHgZr9gYaAxGYohFWN1Pin
DNQ6uNCoTY/dpfozU8G5468uuXaD1VA16bMitI1+Nkt9iL22pqn3Ls399G5sie6s
vH2SdnP9v0+YY3Q6aU8URKPFJFUhChgakvKcFc72iWyW+N9i3PkBwWGG+DU/ATqC
ApHDwrwRYP0W4dW/aacTkKXAUzasmE2waGjceuOJztkZrKCCd1meG2+3JKx3c6Ge
DYJqkrznTo1Ivl2psyu30sNwk/S44ZqNb+H0XuqozxsZRvWkEJ1ZT56GZOh/BMlH
t/mSYmr62EKEekr++oUAXes6nEMG72VoMbqiya+M8HDsLeJGFHB9RL+CPg7LH6Sy
/GWJ0m2RMriU8olBgYlaLsxMceF5FmDl3dum8pb4DDb0x3az7K4+x07KxSwrXFW3
sT9fgxQP9Kq1oPX+4l0OfXm59azoftNjSvfQUMTvLoWCkZIEZd/bLfqyDFqtlicE
DFAaAdOhlmwAdq1ObKb8ZBFrNL7reyPu3mgm9+xnu8D95q2ibqqs0XsWCtmyVZyP
mKQ/KNhIDieX6ZvMDdPNeVLPZQ8x/wyX2KulcVHF85Bb8aw4oGN/jpxALGbHqxAa
N0yZ67Wsiujq5pctLva2TTF58DLIJ9VoF3Jsp1yASczKODqWUFqCQxRfltWXgxAP
hnn/rZYO6iOiHuqmzDK6fHaDIW7w6x1/vciPS1axvL1bOl4Qf05DZLrnfFxURkfP
YpfhYP2YkYQr8EmIpoOcNIvV52rxKnC8BRxjC3KX2P6HzCwEDR5dUZ50W1kZkw/M
GDKBv5MlQMoVqh3Up5Wh274WKFJ64ouqpGWUE7QUUdpqMWz6/93+/EusHZz+v98x
2JRynpp4dN1OAkXHrhiXDm1lRyhTodvVx9ePIq+LaXgdvC7Em/c11DPVoDgvOj17
5/zrztQXLld184bCbwMqCtgTp77iE0GJq/rtcBmZQRIpAkJQHPnK+L9LHPPD0tH5
soyo5ltKTWf2k2KUaeMpOkt5RNtw3RXtPPk8HTf5ECxx5Wn/nF4xRGlNk6S0LDjS
DXszGtUcGTUbMOJ0NpMiBAGGyzYail85ICecsUWrDO+cZuvM8DidzUkylDpH970E
64Ki58o6WMNHDgErZcWz1/6W/Z36b5uAnHKFWi9h0hk7mNMjEd2k+dA09vYplnmI
q7bfVqpBOFqt64eK+jWtxJKRLcGLVXtEjvA5Fivt2fbhT1a2Q98RwBoIqJ5NL0ZJ
kd2oCjj4gpwJEAj03hEkmquvlWvWYTPHbdWM/Hfsrf5OlY7gl2J+ooVtAPdPWQbp
HE6a+CI9m3vC9C2gXFCIz4/sy5/a6ULqK9qam+qJUBp9YdhEVZUDyA2I+9K+ODdU
M6d4UNIkgbaSAgvS8pCgdQqx6iXg1Lcogvyxt4gmttMiwmJiK2bqCqvvpqZO0OiO
vPB3gG/FPCh2RTLWPuxEw9g97jYtyBMvtTI4HiJ711P0TvbnQ8ByYtREfdOQ9SDg
rb+n/QiVYtiRS0ScftDzuyhp0R7kmNTNRIBa57xsbJAzn3eglDScmqj0sVobYwhK
8PIlNd87IhGHZboz+Sey/8/R64GrY85h4a+hKuKPY8XKi0imgulDI9uPfEgVN+o0
6EooDMls9+l/KF5rOM0xcSh02uqE5s/urNLPan3f3QfluMVwZUqBY3OrnYB5Vduy
NbTI6y59vOkK1OtZY3+OggiuRn+M0SZ78FmtogQGSHmxamWRgrp7lrAI+QaA4RaX
mLvWE1Gs8pbvwzUpbO7McUle7b2UzGLAdr5S41mGQsf0gYZvQTjxhen3NGQqqn/X
vH3zzu7aSIO0Bp8aXo6YgtNetjCpoLVcIKpoOHyhp3fZXygrqO8h3zVZFWHC2Ukn
eV1XsoU4eWhIpFMUxMNziqV5UvR0o7pm/p/fKKod9yheCPZ7KhB+jyXMKwy6uSHZ
9UA3DkXdTzLBYAmaneBci8K/AivhoJv6MgfXODrqcTgKL4DVz4+xCZip+t7QXLR4
UXlVbaywFJ6kihs1/JPe2oXENpP8xQNzvAXLJzD+Lkny44hoUON/ZiYGxDp0LRxh
AO7g8fLuT3BdKBtzCCQWFWXC9DvJT0AGtlGlUHfg/ld7wAbhVrIoPhlC8MdEQQUO
9mPlDSyCyVlTwmPk/FE+uwvtQE9xVtyqy4RDZcuUojxdwCSvNn2inv+Soeu+xLlv
jAFip9N9j8uwuIkkqY0TGnkfwPM91jX6qZVjUKI4wMVitVUDa4+VUqsWRmroLCgw
OHkxxnfL3+LflV4F4L6XC+B4yC9GSG98ZjNV0g8QKBryIrsZCUXhCDyqxXBPfskJ
DBIhvh1nUuM+/ZEDS13B1ec+kLcZMhJBGqs8Tg9u8h3c4xUaQD39/75A0zLs7oJf
YfXoYORxz7ddzww/vTnvgoPT9Ncu4ykmSTOk/+gWGTEPwGmWEnRxe/nUpSGft53j
myID6epsyd6GWIZVe/T5PMv9vDaxGw5O44vA0c2f8hGXfY1zGbFRloCj97VFNxrO
S0cRG7rPNtAeVnD5rFWnbfGA8pMCycrKXgBAR3etC6esmOjFNuHto5TerTq5lhPx
A8TH8jP2H2Quh7WR35XFPh5R6KX9EUMrnHtaEjGMhzpp9IDYDMwUaXv9Hf9+ADeX
/O2LdNuNpjGbGPbXMe5y9zf8RMKDH9Vg7gYDLyK/Voisy7ViodJ+UB1Z7+qC4NRy
95ZBWdp4Z2rgLbTkb8Z1ApZn1uN4a4SQ+COGw3RcfQ/jktxxiG+tV3lV2p1xRjr8
vOhsmiT8kNswgFmYUQTwF5SpUEhQOKOm3+p0UMtKrUQaZCDLxjfoLw09bn9PgUvW
6eUSjE5/m8XJV86VFPSII/wROTx94lfQKNIvJFwoPoZqLiaTE2jAqct7dMbwTLV2
AA85gUHW+sHQa/NQCiTBPKWzk1Y6hXhDdM9fXjnzFILCgnlK4qV9CgfDn27LxD5c
JX0evjOXODCYVbhm9jujdHzW9hy/9BAfSBLPei5jYCiuMtUJAnEyjHvHHsqBTkf2
eiz1B9NBDxS7BWoQil6I7TAGUCNSnmS9TSaOoEvfaYVeMUB9vGh6Edc/FxJxai2B
WfA2A+ho6jX/gY3VdF8WzKjO89aim1LU1bqopWyGW8k4GWB2CMEmB/psQJcEO/DC
z2weQU5OtwSLhSb3rF9IuTbXhKLZUIebc0E6rpNM4m5Rc7KPHUPCdgeqPx3WP5QM
nsQ+dg0DhQRlQbA5Eh+XDWhkLJN+3xdcYO1i+frLzVNjD+zKVQKrZVHDPmz0U6vZ
huzA76XqGW4XDqtfKk0yy7DGC08v9OOjo7hbJkLMVlVTX8zaZItgvXYeR08yLv9C
FsTarai4dQZ2hNcbMDPL8uXhp8VDKJVdGwkNuLmLv7y40ELQecy/oreNHbqTmdUr
qOv08f358uG6efrxqua/BG4Rl0q2pRwPmA0ZSvSicinMDisd48zZNZvvsc3HUOPx
PYPigmC0XQVazTVSMwXembsDXG9uGblHGpL1597nvmpHK91dqrjZVmiUjuT0M03x
LdPQS8AMV2DDVPV1wY5006OW3LWdTHW6ta1SHWalJTa0eQjwsK+L0/6LV+YKxVJQ
wQYnleQRXImFykX0TRMJj+GpZcYYG+tIq9SSLXeWkgaKesWZKt9PB1Ez9gnuAIYG
pF6EnseKuzI6UmV1gRbEAyw1ICwuH4naJqSxmOqZxpI/S0qlx25dwWA2e+x9531p
fimaeO3tFwjV8SMUt1qG1lYhZ8qbf/hqdw9u4Jv/ORm2LADZ5d3PAh1biNTJo2ew
ZCr88tn9kwkJFDfQmJEDD4F53UFmWd6znL9efzF7D9jP31X8y/HKcHVdIhsS+2nA
SjeZPFqv3fyqLn0hvJUv81PKOIC9ESrGjZNzA348f2LypoNoxrHkeZ6RMAy84rxA
QXSxwqH4DAQ83oeW5oll4XV6BhAAp90buEWskIlr5A4u9CtQnGQCQYL3ZgBoILvF
SLRnILLK1PTF+CeXvBOM/zUXF0EiyFodldJxJLr+RvcBR6Lp21kRZXwDIXc9jGwd
LVMi54hnOzqJJfO/PpyaaWok9kEHEjjitP4XoNAjrwAjVohx7Kk3Bfis82bvHE0B
vnhrCSpEjBDcZyk7hyS+knlp56U4HkcX/5az59X86Vt8J1PXdtZ0liN7dRvUlBgB
t6RemPwcnqOId4kfN8D4xf3/Df04Ov71QHTt2eJyR4x/o4lZTw9xed9WX+OKMlFl
RVuTeHKv7sJ0JMuYFgGpDK+Dcq8dppKaeP8J0wcVUo0Nlp6lLww4b0G+GPcC9QKo
tvB8gOXxHlgEHUziibkg2YsrAadCX05FLeQzFzVBf8KKsancNrJMy25xv4LnO/xo
dWhDYoFHTNB5Pna0JbsDd2NX3Pb79+9IE3KgwT1gs5ZoNJoiYkF35otnvImxUoza
5exfE7yeOWqdmXr5PJrG3KGT5g6zjYX4wI6P9Z+pAOpzvp/hrm0T60vbZ64R+qQq
XyQLP1NiNJiv6EWUwe+j4tka0qbc/B3qUBNTLl10RBo/lzYeLv5+gbHd7wv0iOiv
GBMyPDm08OIyEDf0vP2aXJIg5Re/OsQSGMbKC+FVu92TT1QnpQ658wV6SUqZ21oZ
da6sW/VV0ZC6aoPPyx5rykzkZQOet291UFLAppzCD0cWZBG4jfDJSoevhDJWnOx2
+ZL2n+9yX5xjWusjDP9/p5dheLrhnKuXINgylozTmpLUzfzFvKlpPihwZIW621aT
mbQYcO9mIn0vDXIG3X9qJ77i4WqkyCDI5UHAZdvuBUG+H0obPXKkwkaHWsT6TM15
bkGjACiMe+0abMnaMVOmlbYpbpjZG1+Tv8Hownuv3qXud2YhDle3Oiv17EVFKfEq
tnEhcI1exsjv2WECJ7xjlthAO6FQQ1R4K19yZ3tdZKsPJuiCpiMoj3eREGuUOFKH
yGr3QOEcrFP+WPidiMNfiPbaN9CwR0e0e4JN0kFHeH8uY3+i7kAnK7BGvNtStqRR
CleZ11m0qCUqPE63dx2u59Ni37agFNa98sk5xU/chG46BbpSKk9wa6TPypJE5fSY
eyDwXB6GrD5Xu1VmFBhJScoNWJQi9Mfh6vuwdYef2C681jdXMP+cisPXrXcvdgMO
JFRNRfUsQEXiTLvyRync5OYwfv8hiAF0RIcDlkFWSeTv+fQjm/uq43VzfGG8sQy2
2ljJ/LlH73q9ZUaZUy/GlUxbpHeYlVr80ceBDOs1kRIcap4oPrEm41vUszAvcvme
d1LMqOf6ZkTXvhcNm+OVq77kP45aqXvvioQlB22UAm6EkFrr0y0nmKKZDjKCUJZ/
ydmBR0qEcYVWJy56YxGNQ58rRuGDW1eTzCuBrPmOwcpX6+XVYhYHkJYVX98jLaJR
MzY5gEWIjYwr8ZhX9l0StxzGkxB77wiXtH7BocdqdtwmV0UNryE19wS2PApeikCF
DpwXZTnzX7w12GgOyorx0hPNU5YtMqf0B5VeC14oYRZfbEMd1Jm0CxhpqTmsXTxa
m8G/dVNUPDuBAG36sDXvYH/3682ovRz15Wc/o969kKg3R5K/hsec0UnQucGc54Dr
jf3GddQJvMnBtW+uqSkpIZ6lRHh2kxu1apuGzzXD1dO3hZPt3J4cteTZND2IHtzs
JFcj6+5VylwaBA0OOtWSy6LKtjslVk3Be5As5EbDIJ+4ZbGvkqDLnra0QFhB/krX
ma1/vC2Y+7L3rHg/tY50+lhlKbzAGRwW9ThYlG5kliWinHXrBaZzieeY/h8vEydL
//QAYoNvZgy63LeKsIcX5lVTBEN/XIhEZzqzPT8RbehIRxMBJDMxLElKZAiwWn5U
kusYC8Q10JXj3smuF4ZSQtk4cLhCsox3ZAHObsF97/8717/YDchp+LxB49M27Ex5
dfTaJsV/m3sDS9RPnZs+LUzfhWyGbtxOXJrAVMAp1puxw8UdOjWFLGbCln3OPS2u
hikE0BEmhyggE7eWBDC+odH3OSGyf0znBGAmDY+RXM+wU0eIIa1Kfys8/tYFnZVf
NSn1vHbxioTBL0VspBAoBvaT/rQs0HpmsTyt6zGtNJ+1kO7zCVh2fvrbyWuPH+2G
qWouTAeO7f4jfk+gwBAsp2FOac4kfdLD7pYxVNAIVNzegNyORFSiIuiFWKSzdAOf
oIi/3V94IMVVzV4hsh9VALtToiv0aFjohd4YW2CU+rsEo36RuGQ1uJZd0k2uDxa7
WrFlyYFOum0KeHgGeHku2zToWf4mU3aMLbGsewgj0oKjBbebA1cc4mEyIg8LSu5I
TDFOvxLf71VddnOK+5wQnRCkq997gf87ngwFqY0dX57XG6fostLMzKJ2momyBiSs
XlsRcyKBKIAllbytqOae7OdztaDWqZTTIBIRGNrNxTi88TPIa+/xAPw2yKyjrIS+
LeUh0d5kIyqMU04LTAnv/GjN+Nwe49Nv46TeCjc5Qqcdoz7CszkkB315tPNj7zNl
ivBoAu58etVhpUvAq/6L9P3K3icW3CQj5dY06Zqhsi18j0LG4jLe8GQLRNjDEPv+
6dnjm/S6+pxdNo/gRjg+SoqBXfFSISjBINkc4SnJ3v/Jppg6wP9dNJhzjVrjFex7
N6wIig9nTDvjFngSKeIzw3NTE3y/pkC6MScFlW6XpmBBnmf7LLui+RWO4E6SW5Qb
twN667BDYWwHn6BFj0GcINNu4FJBpVa72U+gmh71BD1G1XmhIZ4fRS0zwYAa5Xq7
fOD8NM5Vo+LxIckkC1hTdSQQCtkKiqVgYZQJ0dfxzM4zvpeAJsM53/QJcHKEXLl7
O07mZWeYHm5YLqgfZruZO075ad3n1vWZ/+kVBOrvLFrGT62rB4Rt+K+OUmUS9amj
LPD3LWFGkiKMKsrCtxaLL0YFRE8WpQuCm4xdt6TNJTaQb8+IBw0aawplHGSQcH+T
SY7n5zQ/cgOffZdgcGRRGQtBVt8yuL8grWx4o/BX4D4/LRt48+AmSBEA0NphjCwP
8LZp4GjW8lOb4z5VJY7j3C2eVoK4RqF/3jVOfSME11hBbF9JdIkbBolhMsNq8niR
imxu9K3uXOGtej+Wwod9OAyTIELI80pT5FdrzKLrx2X+yYJBBZF15GB7Ij54o77Z
tSO0HNS5sSHDK221HlovDlt9CR7yyGK7W0zJx2YPZZ+buR1dTJi/ZSJj1Xw5mTz3
a0HJU2dZGEzcRfn2ujPWcrU0Iz6MJooRWEcuZPsPiiGvPid0z1sSf+uPPF5SqQeq
OGVh6CYLqiz4WTerdKK5l6t2HScCxzpS7a1mzbx1eFtIr04zZCc/qAXYYTbIzLMg
jDWAk3fCzhVMY0LkTt74wtU6VSm8ZzLEtd2oHX8Jo2IO726Pk+mse0//pgby78tZ
fl+w1O3vurP6K1sFoJC4z6BfHbA7Fx4hSJtry8TGaAMrHAkgkQ7Mu9i941dwBtJF
xkV1FaYRC324PGy9FnU0SaXkpnns6tH272gllD06PUJ2j9n+PFUUmws9jfjioMNL
+uW7d/4QXz6cJOEk49zfi7YSRN1uDzBByxYiGH+rZaMypUub/w+34cGOqqNMwr7j
+OaQnQHk8enXfl1L0wkc5Y8vp0FWyrw+6dQB9S60NEMBvLW8chFyq1kDZMsQrDCX
zSG/ltByDiM+sVFMDe+2VhLUW4w4qxgFh7MqQk+xby32GeH66qxzVT3IPC+pKFdM
jpnp/6Su1zuGHFzFXaierGeLV/ktwYvqm96UmETfHSZRkDlzAiqsq59m2qVl/JV2
Acv/POKN3KYyUQicQzd7Rj/Ck3L65lQf2EYMICgc3lvynaKHw+umegGd5SrNZa0U
p+T7u2gOg28zMiygCnpSZpqYncRFEMhPaYQZRHkIbGFMPb7BbGI16SVPYzn/P/6R
nYXr8gMIfrNB2o74fn5Pwc49WeiJ8u+mIka7JIxK9wyIJP6hnayo7gx9BfkLQ/oj
/czCaXdtOWBvSmAMVahEWGAM7ITuQJ3Kc4roqPtCh6mdigqBMw6kPiaKKx5KDNVo
v/2bCj/XqlPUzmuX5CcrnOhRcQOUlOf3eru6IyUcJRelEUz4SqwgDh8RqjmYcCO8
PNnchgJJ1qarVRq/chY74C9xKRfFiwbZzYIH+kLafMHv+RX0favO8KvIpTdqavcx
bFKAmrjg1M4tzMKiEoX9p6hmFTHgGVPMb3vB03Gqlix+Qd/ZlWmkzr8cPArmC+DH
fqyB/xYYnGYFbi5sww36D/wMlq2d/X6iuIlmLEDqGSU1WhqHQBRW0C7Mo4RCK8m3
jgP87sJRqSOe/Kvl1M7UFZW8iYbpPEafm6bavQraPlKGiRYoizMlVBLfkHmgNV2m
njEOKdLJKQ2mCXPRESJYJS7xiRnbY0SEI1CX6+k1ZFIQTdzIZxWKk7P+aUsSj8gM
xYVQYHQlY54watZuN1y2bysToiQRdqbiN8t/QxKonMQo9cd8GB8aCvTHs1ZHedz9
v87Lj4RB0bMxJUC/UqtBARroTCb1ldoI977UWD9StCEbN4lmT9dJdhlKSz1PAPKD
6EiiUSZFHSE4Vci0W5M34Zf6tXsNGaakA5Cvvpo8Taev4QBGibU0gEoWo3JeABsM
1folmLH7YiOTPo4siyOkHqGt8Pb4LXDRU60pEjHfHHA5HFMPnC1CyAWtxaP5koLz
9S1fyeDqKl8oZBsq8Ln5hZVIJthxXNsoLtH6838PlyVaHNpXY5fiNPCW/BYRRufz
5RBo2BAvZtZpf8I677BXDhZ0jm4sjuuznXbRyg6B6r6E55xSwUfqiJrPofYw/UUV
Aiax/WBM0zgGKUkHZUTEBfwdIY8e2pL65acgWMBALESh7ybG4Os0/OIfn51icX94
UYAiOXFadBts6MUjF9O7JehUqkKSs3jUHXbgwMXrKvzjtQ3Dy07qmzroQxlDEF+8
RGsQhl6zyxRo9RJ/ZaNIuvoYngHS/ASzy7gfIB5IW1ZlJg+7bKNDYN+QopamTzf7
YyzParFrZmPiveU0e48MjfsGwJCQOP7AejlYWiRrHuc48MsvgzrY/8qNszGl0TKH
GfCSP7Au/RsGaDri0W0LBNZwnO7xftlnfdL0KhJ/4cnscoCeJwvXHdkeBOdwwSFC
1dTB1/H8quzXkUXzbDr9rA2w7vVEsNTwY3jA9Ir9YrVGChKzg8xDg5RowcnSBquC
BDx8LRqGh+6oK+iVFdCi1Tqe43iZpPtiI4CqUAlioxfgeQzPIFwwCYmKidaO7yDy
sBOfE3EawnTVGfAc2l2d0m+pgNutnyb4G0dyg9tqO8Ctt+S8HDfHrIlvHZbl1BMW
mCtYoBlT7Bf19xdG+OUj6FfJRJ25+axzLAkFdu524hsaGzqXfnzguaMpcxry8+9N
971XPVaGFCliC9ciHL2y+yFt9D13w0hHPYbslI3Fv6hRy3P9Qu030PjIkmL/ByUI
u6t8kNvqFn+ys0OQlGTdfAHkb5sRevqhUOOk+Y3aKYtOJ/BTgtm1Rw1gkIWUsDtj
K+fCkDNYc14CMBD74pVRcXADDZ/MQCVdWwnwJTC+/HCbDAKMBct8CrPJHkku9SYS
ytddHGfsjQU6QCwW4FeTo3UGjQJn+9DcXjRINrtMhCH3W4OVHQJJxwXydokMQ4uU
dzpWnP4gBgiM5NKOPiRIYK73S9rjj+mYAESpkEqhnGgfxqeU1sdEmHe7qkvYrNXD
fmZXocoHoNg4BJB91ULXHobUTH4pGjot+xGQbpBbcxoMscBoranNQOF7eLHqLFEx
qSRlMWTVNMrPnqR/P/a38x3xTLAH8Nmbr1JyRnfjfvfyruR/J2NUcmhqyKBAZYIX
wCGJ+ZPZjTA1wYNLC6iTlK8o5/KLl1YoGV6mlAm5JcdL45BTlKBGQhgc/XUMAZVt
yuxP1YPkPCunBv9Cp57DHQbk2nMPlL4TmLKMwDhiZ1Qx1ghmG14QgoK+o6aEuVCo
0YnR1MYEHq2V441ZW/BhfDeGOBrn23f5lWYLs5cl3zbIe7YKxTJzPaNKwBZu3fxC
JVJ+FJpjEBbR2LwL63HTWS5wQj0iZyoK0WlQtocRcpaIe50q7JHRUAJrEGmE7vuE
V18WYAmW7sawzZD3f8/GHXgZNhzIa7TEG4LMlqnNF3QC3JEnHNoFG6t4lDY6/dyw
wIfDaWzJ/r30Pfef8I5yO6hxSwUZH7+rVRq7RV/df0LenVZ2SWbpWBNdLvGd/MxN
ryGQ/8S8e3HAuq8PTfOgXimYDZySPSlsWYJJxCI6TuI9Ntml75AcG41hGV7W7WsG
MN5wCWytliOIVbe4abrFqPV/cQXgby3WHS2kfayJEcqa1pz9r3b+sK2fvPmuQdxB
X0BGopq8xopTgQ4gDtWfL8FVV8JUPntq//Xx1PvSOJlZlFNnOPnhF66VqyP8Hvyx
SG7JPgA/mfSkHSILeNkQ1/Gyvpzicp9t43dqQgxqPc3mJR5v3ksUg2pNRYm5R98X
Qqw07PUPT57q4RTcQEAPRZR03Q4wZJFbNH+rdXkcUGB8hpRaa9QahDftFsjjIZuw
YvuAreoaqfxYKQBlQCi9yALE3zLwTJSGYLPWF3DmmNiNuSiVtnV74GuQ4i1gluQB
zI20J2zVkEsW/TJeecZ8cUIOTEp2J/HEHwxh1x4rHuUnWevcc1FGsgNsMc7uvgmU
TWilnbjrZHebLUXnw79/gehxf1yZtdp7R8QvV5VPq78BOtJPDdbdwIfFUtbHwoQS
Pk+EfgHel6Mw9GnzTs1dZd/tU5waoinvPuG4f8+2jwWhztQsWfdOFbWgP/F983OL
+F052hmN79YVmvRsZcVUYMW88tp9O6/lZSDBLHf94rAwWfSmF025jDmtQivmEuTe
vFVXRQmkPGdrw05RczWh5HF3JcNcoiCGqtjY1qA061UvIbgmFf+3+19lhvFtpq5m
1uPi/0X9VjgasJMutivXGSDCxHe+iMahYG7Z59tPmDUxByO3+fWBY70MsvnfrXOl
PuX2SrSAXZkXg8DZBa/5y6P1RK5Oxw/GsMK2MKdNp6WMctmLsPnDYtB6ZzofFyso
BoKSn8ev7UeJ4ggK72zXIZZAZDMlcAf2Gwe8TK6+x6CHQy3unLTEKVoYfwBuJ04k
OG+Fnx72RCt4VfIew3MaA+ng3UvhT1wvqBmR7TM+ug3UyAMxPsVi5QHwzI206R7R
9fJ1d/1CEsRD3sRXEog22uXd91mnhA4OVVgZbZOh/fN269ms+IDZhhwwlfISO6u4
RjI/TOkbUMxhawfbO9k6hIzk2KilZu48UR7U6ArcQ1xF2Jm/WFGIUuufhctr4GPs
xaSwePqRVBQvkJr/ndLgCdIb+7Ds+mYUW5RjLIN5i7qTnrVHc2eXa2294RHxmEMo
4D3PqkS9f347T+ezEuWM0zDsXhmK0KhhZr3wO6UgBXrbmXwQyJMiQo7ZCj9gtoHn
BDwfsH/7kPu3GjfYDZ91+ZPSAO0K06THocNXMt1YdBGH+5Xx3EvVkIauDAX6rBD4
Nym41ApU3xCEgeK5WNywa9eOEEJxnAvENzXD+ikzXXt3d/q5a6oWk87wzUTVpqWp
E9Z1nK/SX6vVhdV4XHWIPdy1gtMXDRy8yiCyeOdTUO28kr9kszRzN5S/oedxHTZK
/XSt73hP8QEzX5B9XVuUYY3ZsxLlZJ1FawyfQrnv0KqdFvEe2dKcBrB9EbsUN0H9
A3i6vXEWPgRC1W7L3GMlUq2h6B1sYMeYXbQobGSb8VcefkBgSfkS4azM/ydxQAPt
KuPRmX0/l0gA2sUBx6sxvOh+6lGvcPnZiL6hXVn/YE3I/QQgg0n7ov9BSq6g3au1
VOwEtqsuIiouTSKS4+n+xx0KDPTSB8z/q7X0HhnX1h7d3g2ZyXPrL9xKbJuJIdhw
SK26y3m6j/plZK2L16/bdu3qNsRXv4wbguUZVv3zrw2bksyZvfgYDz8K6RMuvd2D
wg2J96tQXr55s2zYb0OttF17gD9wi2KTRvXHuDi88MVXMNUtUFcvlIpyBM9d+MG5
PPlNuosFRV9Pkefkwhg9aDKZTCOw0jc1hC6mky6oV5QQMKN3K2jW7IOUDSUNeVxK
8IKUSkrgYM80tg7BlHJaDTNcoB0LwmUO3gdHu6V1Lt/4C3XyrF2PyMZsRxkso8iz
lJMhPoV5bo/s8SdvaLi5illigxjROFVYkF2ffcH6P8bGDllW20g3AyFbbslZGG47
PLJEcoOCNABXI9DIiqnGoPSrhk/RkAHBaoPFNRVmLDavH3JB9scuIyTHBNF1Q4Hl
OfC/zTSoQ+m4PpKqTIDrhI5Twv6Vn6pRTlOBX7XKG62569MQryDAbM3xJt9BbnZM
RyANuFcZNhp+COFUTgazuxDvNdOpwhMtLk4yb/XWVtr5rbaqjNRN+zN6Gh8NhnT8
jPOlNdAakr99uR2w1cVaDqfdTYijxO4pd0kXSTyPDfOqsNZ11wT5IgdivsW3HmCj
F8f2B10zh0MwRmnEq9+mCOKvgbkgAgXfDmXp4ajfRPjrecwRAXlQwkRTTLZYs23Y
KGqv4XOPnGhngUQdOqK6ND7ouLAJIyxpixGFRWyhWOyOk6qD9CUim0xQI8NSK6UW
v+cL2g1eewITj+bqjgXkK4tEk7xZZ0Q2awxbIAvO2sM6eNwNsfsRN/IH5g2BbayL
Qd5PgPa8Dx1Bi18Hk3zB0A/KbpiWZUU/LcD4t0vAJ/EMC9N2mO0OMED2pGt85EDO
WwvkLxzs4A80XPnjNJ16+yxbgUtZ6K5M/AbNny2d3ZSAKQyKoEfmvFaYd4FxaQW1
YHCaKscfrenVY0u8YayNLOOvXrpfP9kZXD995JPlaBtpboF74T4byWjJRqzKidd9
cio4GLWldxjxItyO9+8BBr7d51QNZA0hhRSb9PwPjw/WdgJKdldfUaq3qnjlmyWM
jXFzN/61/0SnnKzSoT/KrElyeStLgSvJaHiIBhLmX0kY5aJKRPYlS26MjyCdLcoF
2Eqnqx/q2opGTpvZZoIu094R44TieWvgWhFX+VariM/574swTbZNLHrqC+PKUB8D
vfAfJBvSkLUh2d3IUDAMmFNZeKu+dl6yonFu2HQRP/jSUAcEDc5yBfrKK8DgpIxG
0TaBRq49zndz+rFfRF1mGsn5dZqLKrPQIh3zyDlpIofbdvMjTBdmuw1eH6xw2BTn
jx5/Fv070my5AC2L7twb9dsv/H630cg6e9nW1gLBI27bM+2okzlKetdnwK0sFEvY
Y5AvOcC9U9g+CHZ9dPxwe+vFXRE2FhUwIW5nUYOQT6c0pVRzqMThfZAPr1G5VfVs
5Je8NLtr8FmxBciKlf+cEpSHVIQMifd1r+z0Ucn8FNf2/n/UsCuB9W2ZFSCmW/Yx
797SOobR/gsC6abNzZ8gH73nkTQyvIOcAF0enWn0JXBhEOP5M3KOr1OqvG4JA1YI
wtgdimdaxW2VO9Yjxx/oBbLPxA62CrOmv9Bc74LlKg6el0etHjJeHh6zTyTeCR//
5fDkP5maM1q27wuORWxcJeO3xIex/CqR1/iTwYqgRn07Kb43O1c2gNt1v+zzqtVS
TQzdyijAmCumj42UQGBWsxQMdA+ozgcOoZl6w0CobdS8xSFfX5IjreKvf2oQq+9K
qamJFlqXDyAe5GRF+0uNzUXKLhHOCQYAPIz9BQqTgvd9gO+kUXuoZhZEpGQrndcg
6/nLk8UdZ4/CychUjUGgrDy+r4Bn7ULoowpmp0a3sRxD5mi8Oe6qT44LusRGilCg
EmfuZcfCXPFrvR68nquQ7xLeJ9thuC4wl61MRU/pu/2xD+3IPnh+8cq271w9j3G6
UdV9zGGcUpvxC4m2ZCagWe7zoAbii0kt3mqRbL4Vj8xpZWkCLvFuqYQA/6lT//o7
uidGfTODGlH1GbmM7c9LHqM+uIr0Su3RmihOvCL0BCvRUIIUVTCrQ3o2dpjeHL6a
obYSJYfc7UaK9BYVms7wmlsuyZcS1nGp8td2gOdbMJkRq1avUX+LN18JnSPmfNgY
XnpQAUQAYvqlw2hC3VQbS5msp7aAnCZQtKExpPXC506/EaXR5u8Oy1bNtHY6VIcI
W5hcmLrkeCq51N8g0XBOH1ah6I4zxX7BuvxVwbkIxPpuKU7FxIXIswWjjWwYBLvM
n5Ufc5gr4X3BKrL4e4tdPTOxlo2gqg4r89TPNjJ0uwQuDwvDaYJQPFzDlM/LurvH
no1dAls11JAeUIB2eEY4lL9VMXX2ocUlIF9BmlPqPxrX7bxsDrM41smW9csNPe+1
XTRJGwnWrqT0C/IZFfqkO/D7PvKe/oexD3U4LPAm4vOvm6pxlq/R4FioN3FVuw8h
cHxFVoGMlEjGM+wzmpPxYc/Zo+q7j3BKv8eBw99ef39KToeiUCjBmmCR3Mt9Y81K
ceUAvOte/4DfaqnlTOdBz+g0KYlxdB/V4I1cVBxiSRG5W1G3DB0JtefzctKiNcbT
z4cdz5BSSjREYPeA4RmKfjLVT6KxRUM1QFuze5Y012KqHClmL9cVAPHLDfya5ozc
smqz1V+625iq/uyGlE6anA==
`pragma protect end_protected
