// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:59 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kn0ZPJXqCcSLkew1YnH4S+A/YjEXewLeGOEm12XJsfbU0sxiTypK0qRWRXoIt0rd
9iZwNptLaBMEIsJoJfQ1b/KoZ0KO34niCl95abQRMQB23WxgT7P22Z8SDwepbaae
nsIiyYhPsLyzYk9bAVtPzBWKQ6P2op66Jlm/eU3H7q4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
f6LrGLPBrIZZD8y3P6N/9v4bU9HQy+hifATZC3pciIN8eiB/rrtl5Mc3pmz3XZW3
7793rtCI3AGP+CpxFqFN0/tItsmtSvilTGbc1caCghq8pqvyUn+zWgnRvNFW+cVQ
szGX0OU1Is+hx2J6H9rebcwEs4EPchTbMtDNbabdVU3HxwLwgKx9DylgzMmWuc73
Lj+LT/VeDHgyJJ5i3RlYo5g+fT8R16lj9bq3cp9HtPmUfYh4BGZN2gpUl34lpYsa
HxOTIsl1pQnmpfWn00Pl3LEmdNv2fegZ/ldbDr1UX3+duM9dmWu67zUwbvFT6Q0D
S3ttXkw4fHyBKfeOP6jZyqK4Mf1mPMlt9I1rkg//INT5ZSUnd4Xb0JiRcLpMU6EU
UTvCzhHLBewzr64jxncj5k98/wST5+B1aGDXQWQnAsYYAly1Qr8UbvDkgvUxzIHa
OAqkx8IAjhIY11lNStmSLG8l1+plirtVKzBZm38RWGqmk+4++OLPESPlZa26t/fd
bxmwqk8M1ZbZx63VWKN9fjD0kH0KcG6jHLA61S45IhQS4LK//S4MmF+8/7MpBAqS
gQ8/l7FRYIJr0nLYgYKof7iGt5SZyn1bAd/Z2kmbF1RLJMZ7pMje79lFMSGyv5t8
ddlXyfm/bR2PX7UKXEiLpf4Dfs15K6NPyOOUCYrviZaBXvL5+jh3dr2ENxJ93A0i
huuVkO3WEhbwKQ4UBvLvTE4GXx9unYx9hLVa0q/wtutZwq7CbazwnZtvHce5/TKL
MM614a3BfmqKp0WKbUgzmYeV8pDp+21qjl7KM6xJD1FrXY3Nb4FS/QHCzB3twekY
Of+yI4FSbVQtfdXBapGgkckHLs1g0LoMlPBG27qw6qw658ALBrC0fy5uKtDAzb/h
5a9AJXDO7v/cGXpXnpEkGk+dRwuOF6OLTMcKRllMKhlJIxriSGzmQk9dtbw9mqHs
EPZhB2M45K/0Fq23hcgoGZayZVqrCFFwiRe6g0L5vKu3nwqKVFgp34wB2YsVFHVP
nN3G6ZJe5191akGZK8r8wJH9Zj810DL678ifShh1AYBk+uhs/DOwGzRjgNb79+Am
Ntrt3gT4cYVmanq7ogpSSUtXPBMC2XwkZbyg1YiI/JK0CkBRZ9HqDc36xSBOLbU9
pSaCj/K1cpcmtkOuDz7Q5yxx1M2o4C9tUaMsdo17NFehGHVL6atwz7JdI/DrNpO9
zCCSyXbOcCH2UuFguRf0iKm1N4KaRgSAMhGc4krvH+eLtfCYRxdnVziXe8HHS45A
6D6AaRyNeVa/bLfR8fZbiotfUmfmO10ffUwjAIT/TBFnuii7ezQ1GkXd5bHgCoz0
T9rtBSizlt/HPfn3pjvhAf6IZRjgODdbcjPpNuSMoY2jbvbTUy9JC9msgdC6n2Ie
XFRB87TswrtVi/oaMzYl8X3/LLlCi0IjqzWt2v2XNldQVYqGcx7ZFJifRIx+YNlO
pVEwpBqvw16ls2Gb2gMHq6hUb+UhxqQQr+De7Egw5cOgrseiX0OEjXBqoI75pkrZ
8RuPgXuuZFNClniz7J5iVpgIO/UeIu8+yxa+EAafg0WNCAXjuyLR/dpbK+t/YuN/
uXq8Uj5jk4XyP56vjSvv30oHdXDkhV9Jd4MOPIjojn9VqawWAjvkDxN8Xu4qgxEZ
fzjVqxrRpLC4CnATSBfOL3trHxDRK7TSWzknQxJ+pwjpEQSzs7jO9vDa3g8Ume1U
jQNg4AB//IQTuUW6rgRhetBTjIsnlOt4V3GI2Eh5UZXQADDSIX4D7upRptSB36xL
Ios7HhW41wgr4wICjntkKpF6ZcMYUuKO+wS4x9L+v9zAdmX5w6CmFU4veGUIC1aG
RX2ZHnU2F8w5vhb8XWmfbpQj2lNBzc7flHGt52XVF29cRhglNyowl75umjvTj6dZ
Wb69I4aVnS4GtQG2UBAefxxePd8xeZxyZ7QjyScQkFztSxDP5BwIcpNKAV0+g0Ea
BUo1aGUYzE/bklNbD0PyvyYaHXFjifZZUGFERpS/ETve0PMLyxrOE6+WUtAC5j1U
gDZnKKNqEQD3wyIGlaU1Vc8I8HiQtJ7cY5zV6k0UzZTrCW4ckPK0j61IoP1Uwyu9
1Jm/XuoAiNqDRJeIu9DehN247AXABm69zmjSiD5mSTfff86cdpjRp3o2Kj32CI43
Q+WuIml7rWP/C3zzHJVAt5GnWCk9/SVv8BfK5LyTS0Yrw+/anhHw9l3NGIJ9mHU8
2ShAxexvlOzbOnnegkmM9p43JPPknn6C9BfmLX1ya9uM7j1gsdC3EXn/tfgFvL/n
f6faGL2RgXqVeo2yuTytgnvPmnT1U2qXndWjf/Ul+jRee5SRvnVw1ry9PWeqvYSf
vUgknTG32QEe3PYMCP7S216xZVahNxqCrtMU32PqPUEPUhJkl/Ji+4x4xSmf5iOW
GDNcVX11q3uTS+TXIW3o4K9s3BGtvOt2XwuDC0rR5OKoL5OxvG8rP6JIPZA/eh/9
ticqlQwmWBS0zPLtK74JAP8yOI418kT+i3Rvamz/F01/1wiJcaFiLLe6/WxSpqb7
mYxNy6QcwMgVtZbkwomnbKPS27qHPIaHPKCbLTYd2/Fw8yLnQY/NUO61Sx6bLkEF
tTQugYP33v6GGWEIGfjWCib5GtOdMcEJK0zazc5nYORhXR4NCXqeaf5m/eq8HP1r
LWhQ06Zbjfof6WzL2/T+R+hN4UAR95qZYT6cwmjB+Q9UG3QEWAhhZIeB0npNzWq/
vRhLeyLSe82a8/5DN+ERq/V+rh8hyaHa4pOLniF4NxfmQU8xJRygc7/8kENlcVAj
IX3SoMlus0PnjcmYJFhTvhDzf4K1VfOb5YxygoL6oR49EtqbuHWqPKJWYmKsN0kV
iCpWfsOjvyQA+Bvt1zwVpt5kKalPSlwwUjkHPrF1gNube1zxT4KXORdZYBugpD73
Neg9mCWGfnJCySPhtyt0JXosd9fmHNHLUW1mOqPGxmqA515bXJMdyBZiB0i/YMYq
7tLLPy+07hfQZ/w4pBqHAT3GANtP0vRs8T1raogIa7b/VVVt+7O75qYz1U0yeAws
QcadzNAh3FCmhYjCn3/zI0fL3bPH78uqf3tdONGHj5UmnPRTlEZvfLuBhS6J3KgI
8I62yl54y7RYfDreiPwX8QbPYCAtxiJ9dXbCi/GXxJxz8UKoofP4ZQ9SdOICFDgW
VcFLooGqOGNf1+JZxwohQuMTchAJvLhGKWPkrOrR3a2+OjkOUUbprFjI8UGtYHPj
qF+9nxW0p0+Ijd4qU6rerP5dL/KAIPqn0eboXN9/sfw3vNA4EBdniigoxdkJC/KZ
fzSMZYp2bD9nuhD6WxJfOYq97f0gdeVk7fWnWhTIM5RerOqor30RuSG5O+E82A+u
E4F4ADXymalT14wubCEecIrEp022RLWWwEaLWhyYepiqRrO2wdR/ISi+bhxUvav/
d1hWt3GEP+nyvU7vKtEoaqlHIU/0EJYHjuOks1bRGKKltYskYTlzTw1FA+3UfHbi
g9sM1Z9mUouijYQMGo1mVgQlPjgUToNgkdfxoJq/IyvRoGreYM4TMcXYLBO1i+n9
4omHIKt8XrDU+xPTB5KRM7uhSYkJn8cp8vuU9XGn5mSxiy6TqfAFy6k2joMafj6w
BKCD3CsHCTXtDBgqAOTDxNs9JjPmB0YLmPHdI2sKJAvVcW1mpylMwL2tS2zFuS7r
9iR4SNLuqY8WEGWtVVtk5WOr5mO4U7emb4q7UE/CyQgoywOGsppOQ7NtsxMHz4hY
Y1zDrfCsnwqPT/L4bw7shFn4rqdd2Am1iE21piM1i2xwRV6EXb9eShf4ggXLmSJR
S0bZ4pbXEIH5ph/5EhEZrJJRBI0O//7dYXRis6GkOlgpqp4+8QAzyctY5rSj96qD
IYnyp+doXJyapWq7R8mMrAGx32h3DqWF3FsKq2PiJo6/cv7CHbvusM+p6sTnHsss
/m4JPvt7XoLaUmPr46b57IFD+whdSuNtbErKfSgPMs6gA7q4HkprXUUWU/x75FUo
ZPEpCSMvFxK7yOmCkKUkCR696NdCfKOBM4aN4J5VkA9lvcmTnag2eyvAI0cOOqqI
dVHIu3QbH1mAASWNv7Zhq0WP/liiEzQOn4Vz/V6MLMxerP1tQGcoZ4Z2k9qMoB0O
fI+qTgkA7/rcn9jpOEYg99IK5p6v0S7VkgT7Dapz9Isd6Op+J+OHJuDsEa0vfCHH
yIAbs63YEevNx78y0f5sYceTvfyTN5tR/oJvlcE9OZ8a+K1AXJK/vd642BEENvZg
0oG7O5bzYQdnw5YcKtkEG/2c0a1Wg8CI4T2wUDoJM2PJ5JzdXSm0SW9SbA0Umrqe
`pragma protect end_protected
