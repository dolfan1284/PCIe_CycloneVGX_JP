// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
S5VCD09NiZ4GOAhYWpULph90gl+R9ZGLU9P4F45EanJqSclDW+PVhuAZM5tfW9L/
y+3plfRDgjBnsq04a27VFBIXshJ5RNiPIJ4gWz+OR2GUEvEOhAvEDlvbZY/NskBD
BzuiLt+vGRNvuy7UHkaoDWBgecpS7QduBoHrdnvqoas=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
xRgHCFG+65+Or26fauEDuHWP6V8AIeS4fyuKnLKV1qK1iGjf5eAzBicwuLdI6HlT
9qS4Ug79RuYNW4M0jHgTSrVTuFDsFPc/9vbiNnhT/8Bgc5H9+8i+ToZm4AKApz0c
2WOXuGYsYyuXlaQXrePQevxftg9EL9gO+UOIHIWK6JP+vePED9YM4NIOvHOWF/bM
vhigi/8Qvxptkbd2XH3j/U4Axd3u9f6YpGtDkrbZweFnWLHRKBV35+xHp7UPM2bR
oEBk75Uqwt6g+NaczdUdEyZIk5T0v+Fv7is7k+FU46pFTnGOIRXsn6cmxi28mIgv
me39rjAF633nmJGgE7AIGVza8QoVMi+ff3wA130UPxYUDanla/DUn03eRBssl6to
t8DK7t1p87TQf4ZPC+AwiQQxRFV9X9oMO61qI162oM0KHL2SycYHKY+/mmBFl8eE
OAU1j36gRysIQk3bnQ/eArzFJahaOMeCGTyJWWY3GKmyKyLez3cJB4qN9Khb6Upp
s0LUtifEh5zS/wlMCDdel/hJIf94u3kx6vqemqPH/Dw0HS5oTDcaJybrxP6nYJ27
4JyYerPp6ncwHX7wSskCAeztP9REQFjxoiyVlWccj4q1V308RExsTUGr0fMmylZC
d+Tgq1Pg2VY5LImhhYlo6Ad/rMtiWRggJt2x+foHUEV6BqWt2fAFHFHLVMNZY17y
sQgfSwsK0OhQVT5v5oDV80trlPNw66P9nCdQ0TW/sRyHjVfkScEGsmx8GsZavib4
51VH50cn0hXPWecBGLpJWv5efkhbPEJjhC5V7tlrOGzBkO6USn013XmTAtizlIdj
0IRlUu+bzaoeW35CSkYtM/3o9/acq3B5A7LIKbIzIiW0q2jKzMcC245SipUpScqk
XeDtG7pZL5OLVx0b51j9WXghf/uyu/4pAaius9OAVLipOy0Mh8Lal5W6jXfiaRt9
EbJgYDYdmBNJ3l+qeU+9TTYZyIUTsWGaJtS1j3KeptI+dm3IL/9BCORVbOyro7Hd
W/kvM6wvPH+JN1gxy2TqCnByQ1SDOenxk8GPJ7D3BF5gqsWANibuZYuQ8U5Cnrl7
Nq85dfO2ouh/cFTWm+8NJVPAgRSFDBQw/ojIz7w7stEKi+tBnvDcflH4pOHvtx7h
pz6p7ayvqXeDneifW8G/JaeNKYgJD6rJUUGmYSo6cheel6irFL85W7WjBspCWtYg
gYOAd6ZV8+kWQNSACDBFgcTMX9Hd9haKO1mhs0QkY9HZunSvnKAXMVydY6RwgqoU
iJuHsyWmwvVz2A7DR5YUEgUn9rHBT7zJVKyL8u6q87emAt7gyCCRgXinorYcA1ar
ZsIlJ6OZeOebsPigskcFwzeCy/ypYPvNyh6b59AYpMcUYosy5UQagY3a/Nk/tf9P
8PymN7GNgkSXL/0CwEre6t/SLVVaw7OUUS6ACvZU2B8N3ZxlXqO7VDtwfkD4DSCY
GBFd8VlCJGTfhiaITho4nSCrZ3goDvwv9MPm4auXAL7+ikec+7qDfJFkprngMpx4
dQFqa7iCr8K4yfRcs7Un9mxKO2mYsoz82S8kJB6Pb8lqKdoSvtFM3rBuzgs4UjSr
bjQ9zxAWdFwY1v7MxptAYlm/l3/T+DAmo9dJO1L7iyOWs986OwyHbyaQFQUwHbLi
CitzurjjjPUX76nwEhOQ991VcmWoOBYGkKzP7Jt39lqmkpxhEqB2AT+CL+5j+362
D9MIxjOs5EgID9JyFaGsbHBoQD+qonDqpjGp/zmQT6peJbtR0YeyqFG96VY8VPW/
gKJtw0I3WXTQuttNP3yHfqSB+zjyuZ346CHMoSIBPFJPajV0jCaV3dCJwegJggi7
8FAX1PiBMM486ar6u1z8XYpEYKZpewhLsjgl2my8m6C7tU1bDOdua4tlBjxfuLHQ
5jmj2UxeTIS5alQBHL2Kyw0ds63QZjtO/bWzX0bpa6VeqokY4vnNvPdLclXdmAbh
wP8dfvZYrQMAdxw+lSdLuLxOwEeW6hR8essWnHf7EU0+u0y4NHVn0GUabRUqprjV
od0vjDJX0Ot+Emu4c3o/CuRogxIP7HYTolLPAtsTLv+agTkW16YqgWQClPU+z4q8
JdWdds0XniLrBp6AnqmVJuKc+21peIBAKE1f6AwX4caVIfgsr2J+Arc5Y4I1TsVE
+ty+U3YeSyJoz6FyQcDpq4BRk4H4EGMS5BMVpGOWq7stZKeEcYfrXnhp5zYs9WJv
osfzCUXIFp6Dt7d5Igj64Fge9u0135x9+zoo6jl125GiT9HhB8t/zLrPkKXSzVR3
6yIKNDZugrv2iYj098G3mrZjGIauyjJLHHwuNM68eJ2PqhNEODiB7jHVqVuiI6fj
uuhpG0BkKbes2xpjyLaHfBfH5VQrWOZKh357bawLcYBY2iOVs8kVpPTG6Jaf+L8k
hIg7fPbVj7Om1kg093zhqmgLODsAJ5Te1wPGZ03CnIVC2nbdCOEHmGF1GSc/gX2k
t34G3jaLGM+4ClR4jDK059yIFuX85DusUOVGaTZ9uzs1rCat7INfpM7MiKvnB6ra
/EpU05Zml/5AaHgVqzoM2k7KajBX62/w8jHGnv36k0w1+Y8CVAXPgqcsULwmk7Hh
PaMmFeG2fKIJNot1nYaito9JzPIe2EbsFfeArBl3le3DhrMLMKIhqvqwMJ+pNdxD
mP3pc6ERaQY0Qqw8qr+Wzq5GoQPHHlP1lABN2uvqeKJR1RQCMn64lhdXJuJHsu41
7RIH4iy5aGlX/8BBGOQPfdzunTCZe/EQof+crhXJdp/gbRgWPL5OZ1tLNIFAPEVC
8Faz7VZdQFcvG7VstC3yzIVCGJhsB1bQWTuDURcK2ewY2aiTAeTOJ1nOvauxAu34
2oRchWMy6HOcx/Js4WGT/EIhVlWN+HjI5mtE/G4zRUDPKaqtWJeFEHJXSoYV36kY
TcGb8Zbx0fZaGyRbvQ5Ouu+K1vmD5/FoA6q7rLUfMTV8twaHtpQY7ts1C59TkFxe
XZxAuziCo4nQr2fStYZoS3tyM3HkcdwkzF1XLnuF4hNWhZFTZXjKzpbVDto1s0DH
4G4vYoOJ7Eg9FNQENe1x3+yLrCe1QQ6fmKFHh08n2TFa0Jhs/kUiZTe8a7bqvz4g
TsrLFtCtRH4RD/31wVJ0v0q5AtOfXqvQhAYZmj4YO/X/QdQNJdRuWvKrQuIbAr7E
/fN50gM0H1Gqm4dveNUNz/5JBir3rPHugvFrHPGm5zdxYiCZJJd8TPns1j7OHXDU
8uNpTJCaksR8Q9xSgtG25g+rUvMwQQ51tpDFMtvD+QZljZJImFbpF4kg+PUQcfcd
wbms49tZrZScNdx23VsnJwGGerLwbLZXR2efPDQONcS3vU6cDy4LApCDP45rrcEu
aZP5i7HsatKjFCxIiCmGgumxciPLiwag2zXELdiZ5MQ9LcO6TVDVIUWiIbc1DigG
VhqYEaD/VZnZpZwuOcsmqpLVV8LPXCuaa6eJJU6lP8Kz76ze3byCwl5r01kSc4Ps
cTqWCBi6zLOhUJVhb+5YVcD7ilxWwg7gv+y+7GF8uZyGuXDcWHdFvF7bBe7Zmle8
+RlXCYochPp6nvn4JpkFIZAG5PL06BFi/LmS78WOmbIK/mDvfhWu6KPGEMrRggud
pmywwmvnE8oo1R1qq4tcRvvKG5jvRPfJFBTqJHVTwYbdgRrwmP9WMDNMgkMV8I1K
NE/cKw8BWnbuGu9Wq3YZK4LE8RdiasJ/DlvUje1oAsjrnGtpfFVO7o8hOU1tZN4N
zr/2iwziU36LVfA+Yq2M501SrIOO741ASYQ5r+Vj+1bLC7vpZzHdJUspkj1H+SgV
gQju6M96WpXtfLHK3weqHuBCodIk2jycxHHS1Q8P07JgM+urHzyF+JGDkjJ4W2J7
Jet1gjqBP7Z119m9gSYySQfccQwqT6Jxl6boh5AF1Mu1wrp6rdHMxpLTSnlJXjwX
pYT28+U/ddJlpAzdpEfzDyRQnrPJ8SEXSJ1mOxyutyt2JR+Z4V9hDbQKJ14XpRsg
0ieDPWKGPe/HuwqJaRApEouJI3xKQnfSU1gp7zCJqwI/1zfZStDx1dHoCma0KM6l
RxpknzlywbkMMTSBL3VavPRJ9+TVoF4c2nCtpx8LdIxakxgz2CYaWzONlMnsU31t
PWIWk/+5Aiivzjwf59MH1ECx+U9qA3mtAB4TmvXtmIuxICwpJslkBozH9SED6MZj
2EwEVVO5fAroWbLe6OCDtxxU+e97Bv6MqKNw6cno4NypS4QK0m1I63+gkL/dMupe
rn0RlpxD71OxIvNBVVo/dza4wfSAA8KIE5LUbara07JEmWI6Yd2onxwuviOnPnV1
PmmcQHybcz+dDx6XfiLei0zaX9l1oW04HX7TScnSQcvucfJuJUgUYOKbuXUnwyPx
HbtrhGvqC2o78+UDjkGjhuVCot5gyC6LSPa2O7S5+xH4+byby1HjK9dd3nN+4e31
uzVzCQVSEruP/PiC18WluxEk/NIY0Dyc6FxNTSYD9dLj4MLhAZaeE+hWz84cWRA8
vX/kUW8k2445xk7kErJCEMUC9673GkYRqxZMTe/bV4fAN9eHcfh+CF8/wF9gXTEf
URDTK3kJWJPPmgkNiIqEJlPsoEMeAAmkIRXo7wmmBy3y/Z99KZUPdox0fR0BWzEE
1h/nPi68MK3hGHwECVoSzZAKhSsq6FAosf08iUd9DhUXH0z3FVZiay/wSi1bXtKj
GBtHWna2R4paI9BfldRscq0DSuBARFbrP7wiM6hcW7Zv/x8nRXO/2gHpkgWD6cPH
ge9U3599J/kYdw/9FIrSPTfHqQcm6AiwI0FuxW21fLksswGFKEreqagaVFVJxpPO
ZBWbC3InUwxT4XrN1DBJCQ8DJ7xd7D+JvfEeTOH0XbSpeOAtT49+tGvoaMjO/Npj
sIGGzcM0AzbNBehfRMlJ3kbt6omfKAe7z5akUwCqyja3uhnWxSf+DNrMXLtsldjr
tMXdIufJsuNtSZOIi38Pmqko7lRxZLutDdK8pNqqMXEMhJEARRnHbDW48QM5j4OH
iKkXeYxkvRa4+fJ2RLJifn+j1dzlSz+eyqYPLE4ctmZRLSOSP6QRgA+XI2gOHM05
TpgdTwcUXL3pQzUYiqNWV8gOxw/4IFAxMua09THl2b266d7aU8qwAQGZLBH9g7Sx
mYUMnymlaPRgDS691smRz7WrZldmP3ui3NdVVJBF5dEK3kblOEjvWo60v8qvM6Vo
sChDYDzxFqXSHZJ3SKTfcqdqHIEIsHEKT3a4PB0GKonougmaIyA+VEUNYGYmy++1
ELXK3BFCXRvZE3EOYiGvtwKS665IcUM21vOeGvSjHZUyZXf8GGUvE0LbrG6TtRrN
Vvg+S1kc+vsnJDoFKGBuFaTml7EhijnjIsKcQHXik2WYqBBvOH4/fjt4lCTyw9+x
ilMAfJbe+qr8imiBfF+9xPFn5sSEq20uWiS6c2S30rgBXJ35VElnXndGmu+MAvAP
HrHc829o7hiEphGcq8aoQOgqE9eoitc0uLXgPDRzkhSPOgV0I+QJ2ifquaZCkTNA
Rd8b/ZhmnIC03xHsXuNehcYhihWvsHG+KD4QQ9FgCotJf9G/KtbMJi0BAOW4K8Wd
3WVUL6e1AStyPyfi9Y+FsbEIQbZNFYRm9XY4N018DgXCfHIrJbJP5VeG7ouzs9HY
26oubcjA2a06SxQVLex2tGFPWpkgbKp0bLcJQ+3xeqPKf9p/dB8Q8ugdpXzW6R1A
OB9uFdRRNjdebV+NLYaLzqVUn/Cv2PufbYxDpYRyCPWJZULIWi34yiqZDapGdSKY
9QYCrJKch3V0X0BMGWavXwcev8uYfclEB93285X6EQod4M1Pu+2ztiWLnHJERgBo
ogfLgdieUh+Oz1mDS9BgRluxM+2mVGU1N8DhLW85az6B79OjAaqYUjKCEuaTIyxQ
0bCExXJYz3lfTEgxhC56wSn2MlDxpWYY6EzyRpHsXaB1oDyN+06MNyAH47NDt0Bb
zciRQ8OA4aFI99B5r/pz3PWi4uBbxH23I96Oy4v2QVq9cvI0bKb4ejA+miRgq3k5
kTpWPRuvw04nWud7M5v3On5+irXc4TsmuH43gRnUbWz5RsY30UQvLep4yqQcf85D
oJzhPlv6O7JxgGNvO0Q3nB4MFu8YgsXO2uKuakjD3i9b7sEE9h67tYa4VWiYIcJH
JC2YxJNchNW8pc6GEMlUsZvhpgZ7tS9rJRrHqmCaot4m+1YeCnWqOekRfVTJB4bE
BK5O2f+9c9Nxc+Fqq7uL5wznVhmEisO0jvJ1hMedc0pMaXVc3wl+RVcrrg4gjPbt
CHiStrC0iG1Zg7SFv3FLHsEiGZdxU/kMkrhsRfLbOW0z18jDPWUc+KftVky+Hz85
3rv8VyX0Rg0eqe4TNs2nfSrAhjFah2LkKhUBQTQeGkLZwaJnTy2iqeHeuG62DOUL
ExF517bIjOJd36eybFcb9oAXnt9tKptpu9dhWmV50bURzLtD3qQre5Ehjxuj26B+
xkc1+9RFOwy1WyEr1UImgFf6tr/sYhlMffa8RRXWPEQKNKXoio202gW6SWvbBlM7
KwOZZ3KtbMO53i+wXLJqfXyfAGNqtHYzpZ7o6tgzOvNpIGlLfXwiqZGCkAN5jCQ5
03ViBYxbQCtwckW8eyVdjo0sSxwIf9Bn+0pireEy6VBVQ0+1ifisg81qxw923XXY
ywlNkOf+anpHiCVxHDZhrVB2iGOJJxs3kN8akurun/oMK6ZebgTnU7t5hHArZdgi
e6db65bLNwX3ZCSlwWvFbJQLKmfqvy2xajgdf8BjmOtCNlvK7D8BLYNxA168feF5
LdJSVbO87Rs7Xw8JjpMKa3QzZiz5sdSFLhh+vxD04LuJY2AwQJofFUrtJ/FL0LAi
NzdZ+ARl/baW1hxjSxi/IJzmb0BVBmc/xQeCmxcvoS9XDqfCjDphG2VQKA11PUDk
Bgk0Yr9JHF6Aa5RW0CWqyRNMXDTCswtME8iyn6JKm5mQD61ROLk9+dtXNw2pyNim
hRFESmPnJsOPm3n4jVOyzr1enCIA9Dcz+3ywo30S6thE16aI66j/v9UfoVl5FVyK
nRVDoQLePR0vaSP/+Zuf9A8xMKMbg08bY9Psg0UCQkASH/RZuZd5RXQr1JVuO4XK
2ZLsAWZzdHKJYYTAog7MKUfQ7wYc6fm9/qYWHTglI7qut3n6/1iG8mWtwNmObWt+
mRqaquNvnzh/J4eBxgr0FKcl3VNgLhZP+N4JxVNcjHQve0/hYp028NHX2oIZ6Ugn
9zm3x4C7fwYiLvFC/bCZ1xYjeUT70kG+SHD1wPcPnp1IBEypXkGJEUDN3FZ1XSNf
/pFlJO5oDPEhFPo7w2ViV6efJCybWLgI24nOQIJ1nmzdiPrUxPsM+dAsjYDRdbll
QyHvhNrARj2eEyefFWlxyw==
`pragma protect end_protected
