// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:06 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jX4v3SbtMgpgOIFtQalS04p0VrDF5T99a0Ho+f/+nFNGAiVRJVyo6QHfZUJ2BzHQ
AhUfakl8HtxJTHe3EJ9DU+1w2ImO34O1vUXZ9RchS/ruohYt9+5KDABhn4CZcs40
Fg/I1YZ2klPreE4lVwxUH9x2k1pE0qhtU0pKj0klVRg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8320)
cZEIcxMpsk26/YehlA8hFDlTLp+UmScgdh9GRT/kp/IsyTUssS+drbn7WWJT4Zot
muWKCBjZY0ebmKcKNClI0pSIVS8ajb4eXdwsqvlEMJMGNCLYlM02QrOedjBrn58b
USVABwd848Z73PJ2tHn3Q2ruaduQmjqPYNDpyp5aN78I2QJIfuD6ns7OISSy1i8F
OnIiko1ogIxGwS6erf2uLL+saNNKDTW3nIa2p1Qb4u6Eh0WaW94mP67GwXRagYf4
7m8LRRltEv9xxiiwMvqtsEBD2jiRFJTLJ3DV59Ah3sBksbtKFCuoslO5m2rGUv7Y
Yha84YMLObZpnLjxcKb202ti2YMOJauVV8WNUQVEgJQTFXEpIVIEPfaAVw1PVJiW
ynW5OFmBUXjGQLYYxCV5VQ6oZX6gYj3+aEcB2iDUsHbtnPgm7n6oj35aKoGoUku4
TowzMuBmORN0wFjZ+/2d5EP1dTO/HVO80fMbTD4Osu8jR6aT+ltGZnNbj1dvmQz+
MQlIjy2GF9VXZMbhR1MY9AOnvMc+0PwbKERp68JoOFSY0zj6Nyw2Dd8ufk3cG08U
L6dmw4Zfwv9NZMSQ0WCGl52lCiV0PQH7JOc1Ie3tGHVvnd5192dE2w27E6cEBLJQ
69Vn5w9iGoGOo/+HKCF4lYG4WxEfqMg84XfBdar8HFm+sW8gPDtslaJjULdxxqn7
FMiTP5vSp7+sMPZibSf/c8oQ5/ExwHo6BKtPm0u9aSF6NdOYLR+A5lUMF0j9esX9
bTqvJ18DnLxck+TdI+YAcCG43jKWecfonEGFJifDBiBhm/ba/QPOamleb2uL+9oF
kLudYPfrjkr4xWPKxjmO45yeucmRs1aAvaAZ56HesFNzI2UqbhmUydElz2wj/S1F
8Y6/xCV4cAi5dotBQsBFGFUvuaEKedLkl36ELz6UJVe9fA4Z7MSQPV5yvH9E33Ir
suYO6hZxS2bQZRebIWbTAvNK8gb2lgQX28VoV5aFydnBH96lXfVBn75e+3Fapa5h
EDbrKERgJ5rsPO4clCZg1AGM9KTlBvjaP5g3JsLPd8aDSErGcHeUGUp4z5ddhCPX
IipRRFTETM/Te3G0BWlFD+AlO/h5SzZaVHFF0s7AF3CVJO/4648c8tZ6pr6F/mxD
2JZcwcMoNxSAEf4UrB3N5rNN9TKIfsfZNuI9eCJq061okXiKM4iLcChZ8DoY05Iv
3yRq+WQEvlLBzUJM4uG4m/MUGHxTZiEXEuSY3cOWZjtBawx7BuMYCYwm3XoSpo/Y
huAIhLDIZ/Q6OM/3sAehoeOCLI/NDSRjqCIUdv7G+QcgulloTdFDBBDhdpoBAsYj
IgTR6OjVa0Emu60MY+B4OR0EStdFEXI5sy45yA3XV9/M1Lyur8FI2X+9xpzjJsYm
85J8mHk12+u+0abC0kmS6rddh5pVXRlMzvgSGYcwZIzCkFXYvziPHiJOIEEI/lV/
pOzpL2SBzL8kUeQt4NQxSpT1b7krkqKEYwyYLT+Aut5EnUhe8jb6V43keErZ0Re2
p5zYKJ17+HoPGa7SSzOoh+2lhO6eXShuINljerulcRpGcxF6Ax4mtGa7wk5A+yjk
j3GKhENoKcz4wXs+OxFZYNMUBxZX8GBdGm9uUTi0A7r0gLwyz1Q59EMzCO36j+db
5LoRUbrg1ogk8vWGXt27QDSzAAp2tLVXNIB+bMwJZ+NTLiu8y7Xuf3qPTAh5SooR
zaBGFym2Hg1JtDEiERfQIisFBg0AHjV6Hmir0lMAXXwACKoPTimV5Ihhbe1Yxaan
A5cCQAJXqYP79DtaZm7aSn4TvSwBV3UWcgrrR4VWAr5Kj05CKL02VkrQ+Gl3yjy9
LQMuwc3QpPS7bIWOAwOJ0rvk/t8EsEwrbmVBMMb2eIgtahX2talNhHMf4yj05kQg
tqLcp4xK6PVYUh/Bbj4SwWNRfUTtKrTF/VbHbIcrglKn4dyGhT6iYxPZwy1eV/lk
KyS9JnMnH6unBGyL14HvJ99bLD3O6/NjC7Y5cN1fZ6pAJWa2KcH7T/g0829+Zfj9
Gq7C5vir73OSTTu6sB8533fwFplX6IKvO1/nYyyxjgfVn0yk5Q6JmQ3adlDWCtiF
u2qSf8sFwqb4e4SkBfMqC2WtRQ3uQEm+LJhP3UhtiV+w3zVMPuaKCRmXDxXMn1bM
MKpeeOXm/gHgwRPOxQogsyFqIqdPAuF5oXSGJZ5wLNBgsAASHkUadl0TNFpqCa0k
gEzpB81hRiieOmhh/+wLLM7nwgXNjciH6ifi2A6dSM+tOHaEVJrClqxdxKhkJzzA
ItNbhtBQylwkylUp93PM+EtrCKG8aT4VQwmL3cuPO2RUa9BT2hvs5qz0mmfKCOLn
CI2klOP91e98rajcFKZKOnV4ecPEaq92F1HxSWGTgQen6w9TEbpBL+CQTzHDzrPv
MQnwBQQNuhcHgEl9hD+cg8r7ZN3JxUG7/m9RKToHZX8CrpxPkKyIxwkuRe+mm34A
Li8l6aQdRNFaQS89UQt1HM1dnWgmWVsyWG6pKIaqDsLKECpcjlNjXmFhmm3kSO3k
OVnAcQEGSMkpeXqrQ8GseLyABKpM42pyq4x3MgIiCSnpjsOE1eYp+LCftxfh2pNB
2hBuBJ1Zf0zZ4wM5NcpE2gusKnq8l4xrGCLW31lBrtl6xYq45HjdZseMqtmS5PnU
h8/GK8dobRkwvYVucugefr7s7vc1f569DV3ZLP/q2HgR5HucSHYVPvLmEoIDhFQu
V8zOM8raTZlTt2Fsto+bYNiLhkp4/hPSZnZHxBeQkrwA9GItzlmqIRB0SC9eqvH2
t+81+0YOqJnjPQ1T9H8OMdtcfl96A5fCMDwD/oZJ1HigJWTlfnvqdNDV3YgAhwV1
sbt2BC0MOGnOO4SUd4H5WaCecz6/BoUZtiWHxGN9WM0NvxTkxjOEoUzhiUWq5OjT
mFLH/WkFTPMmiaz1EjoHZ9ajPLA78KTdcLoPCjWtG7wuFps7qlk+WvfaIHiYKS26
8n0qmpQL+RbrYp1/sCeUdPpvB0JcfaXGcggX4mxRXjLdkpojMLQ/EsWIBdOQJ97J
SEcEmqByvjqjH3mhE8IBD76lHEY/1ofgG5Re+3vkMYPqSVkSbchDMwYs/GA15M6Y
AUAUWX8AvaYEDy0h5/UHCoXx++1gjz1n3R1Cd27SOlyLh2zRbAKVfsKzfsAO2KYH
nWz+5ejRFHGHoSAUpqtz/YHmI80VtDTYA5oTHPwLYcqCgJ/1hCetAEltll0KDhyJ
F6Uxja4PZLLBGn69tRUetOnfRitWrkMuod9yTZoYURlQVaHSFQe3aXIkF2lmYk8C
WLKc5F3fK5at2MKBVBpQXyajcDZoXK5mJQbPBoagWTj+x4Lfl1y5unXQKOWlP3ee
uBH5Ga3ERNU31Y4eXoeMx+vjwGdc2s8QodsGYcyQ/u31VRhS+/kmMYOkmADQod/E
nDA7/dnQ2yxlk/JgwFqoyqiGV9xFy8rtmzNSVdnQU8TYNcG2aSUhKMwnDtTCMYdv
qxxEFXl6vwoZWsIfkJt8sTzEKXlwkIhKXojDR3P3JUE01VokCez1D9L1Xa6lHysg
oOjovWRKt4eVR0RvJBVW38Va3PpNvXgzUtHFmvb/5qr4ac4G7lWbxRm8JlqdDcPz
U36apomM/XBYjqBOYA1WmnCEPADKUeya7evPcd58p55yYfkLxZs5IQEchDjJq+Nw
DMcQ5mKNY4GUW+xdqDKliVJCKVlo8o2chlDG4OjIIPafIuEuI9/XVpgTp5oZ4AX7
ecPSX4MGp1b0vHef85otC2iIejI6grTvwGAOdQ2bA1VzSV0razb+W6mG7goS2801
Wn6D0JUKdwyRmC3DmuYq/vNiQVr0zwjE5VhOSs1vVzu52hpymH3w3nYSIn2toQNi
SQIha/+H1D4/H5tr7/LnPdqI9HoNNKYiPtETmzi6TLsIBdDPitFIJBtCPnkHjvwa
3snB659eAWCrWLKkKrQfeLCyZd/gqXVijvXf5CagpGmpB9EsEGyIIUf6kVEkEhOo
mQKrxe2hk97gqBcNGXqG6igaDT+Rdif3wKRqo3tCgCZ9EqZUhQT2AZMP6e+jNBqc
SelZDYGEyw5tROxVH6YPoLbQMkCEPUCrY4w2NMDwW7DtVc+U6nzClSkH61K2MS+S
qwL4zoHnnDKOmFl7GhadwbzhtdYWC9p0xwBBP2LHrqwz9CVzW4vNoUSkWlu8XYJz
Zr1eoRh13twYbwZ7UAR2S01HFuJvvfg67DE5uf0Q6YP81wP1KrkJCZ2bbPSDWc6g
Z/HK24ZLF8fyt/L6Iz6MfLe/J5e/BUygMIDCXjRcC27uUu3BUAfGlrx7kkBEUyiJ
iOlgqsizFn473WyF96zLgDWV0kFouUj/JKlB7+S+4+UItcR4letCSNkIGty4kTeQ
Iu2aMVf3J3cIsrFilWoWcfZmCzaPxkYFEytRRFzksQ15fMMjW1DIXifDx7cuod5w
Ssg/n0PBft6/eFvGxwj6TH7EqR9gpPejbWvdzdFXvqrYgOr3rYz+QkzDtDuQ/vx7
yGXoVmxYOJO8eJhUbNquzJ8Hz/WX32kZNQndmx0VVbnaO9rfVKAO66bkNHX89g+3
Rc4Zo/JjuO+em3nWRoGRmB9muwtifJ/e+b6UMtrAkC+Z81mBvEk0iRBV0nygrmXt
VQz4x8wMHgkAlMUJE/e5dpzGU8LUQx0GSHwcRRv3nD6ws8rWuJEXxKnVc95uXpdZ
u2d3XhO2MdtZ8p4ZD+Ffd+gcMAGd3YSsvyWqhWrOuZiuaBoICHBKQfUHyvC/oXlZ
HEhhgIXweSQggsCVws310FsvU8PuhMJDfi1WDIEFG+Fh/lvUefUTEvwn9FsMj1iS
ZBf6rrOXbZLujCVtDZs+bX2eaefKt14gU1nOOI9vawleXBxeO+ApZ382MgkCmbo5
Ev7H9+xCQ6bW8ZhT5IpsNK6ZvmQbxsOqSe8EawFKJqIPHPqNOV+sbuJj/9lu3zaH
ojmVMAji7kVsoFWDurja8bLC85oc1QD4uRVdQNlNiPSynwIHv7pWvp7ssCuQOfZ1
exICvMnRzuT7lVrVhD2cd6DL+dpSv0imnZmOOiXP/2Ab7ZY3sCWRpqgfDZ+NdcpS
7FjqeFID0TIVFlvwm66DvsS5folqq0KYVFOZfQfKN2VBWVjgjuIkYZUfgCF33MU5
wyz68f2/VOrVQcAYiEePjyRaLKKE43toSRJA5gQRyr5UGZu/+ghitaiw+Srz4SY/
sDi+rhrKNZEWg0aXfPgc/dIPhl5cl3rzWhKbrkuEbDNYdno6obRYCSEF60TZZnrn
VVS6ht8yeZ5dL2lTeFyzAkaYbyyF8y16tRdXprKhmA+E4AVLqvNmpyJAxIJc1F1v
37hQPpo10XdhNgxJgBqoUhGi8PkeYHaN6tMdw4czQAKK5G6QzGGMlvN1TRabo1dK
/p9kiPcRGet2n5wcnY1sumFDTJZ3MVRQaT2lQ+tHdX2UQfUty+dYibn18NjBnF5G
HfI/98NVydBWgq8fak/5IhO8o4ST2NlUaFvJmSXMgd3uNA6m8y1D4zLRPlogkDJz
lkYjfAxBdJ4J1NIt0rJ2q9JuI06tUzB2sFI13uW5Y60WBa7mxOOWKOs0/Fn8hskl
OJsIMhU6VZ7yVwIvldsVW9Bfbkcq0AB95ycTsU3zJpxVOIHwRSkDmYFaLO2es+v/
Qs9AErKozPwLj4p4/anfronoFt6iiuNu+FFzaLpfV5A1BwhaF0hqFA/QN1esl6hn
ZNz8IYffYWrtpnwLcx8XGVJkMBXohdW6HLRH4pZ1/T8cTm916WnxRkggXpf1/Ssp
HBdRNMiGy0oM/KuO2bVNqLKxEavebXL9CVtRIbdSbAS6BZt+zeep7nq5oPBrbhC+
Pd+M82Z6hkwKgMdT8afJG7RrSSNzC8hjkFz0c7v92Z4Oo4DC7tH+Cvrhn1gKhLcR
sZohdTQ9zQQPgsMjvq4+/TPFQ1z3O+M4o8UF2NTcrdqbK1PlPZg5M5vP3iRAhWIw
yDOpEsLtxurZCSRM+jcJr9e65N+zVg3gP/5LlEHz1nNXTRZJQDn1izPJZYKZxuQK
KE/nSuT+J4Wy0ApFl7lhwbPkWJo5zuCIkI57kxMLzWODX2bjSh7ZH4VPDTk5Hvz0
X0ETdXJv+2PReRzD4lQIDjPcpKzlu0bPaC9RE3i+iGJIZbr0JyUUcy7a57UkeKiC
JTf2urPrSzWN7eVrweaAIbsOQOwetVpzaAUW83mKJ+DkPc2R+Mg6rON99ERwGSTd
QLAqPu4l+JpJpTge7uxhmChpptmXs44ANecABl6OaHvPy9vmTsnFg5XjBbLHoCbk
Z/4aZjy0lsCeljVBI5Omu9odQAts75CFH1fFC5G96GDitZinxCfmSvyzDe7AoNvO
DFuSjEdiz65ZiQeVLGEFVeOBJ8rJRWbbufkzHA9OMCMt0mC/UyMKK3T3yz0g0x4G
Q790IcQdsBeG19Lm7w14sAPaQj/qh24t2B+aLbNDy8E9v/A8FoRaU7Ou8hEC827H
NO98vdFkitFEOfLymYUgI0TWumqxyQ4+2Ra0pCfXvn0BPR6X58FJaxvT5XaAVrY5
qkF/bR39Vit3/fHFy7byIxEx3EDK5bCuiHp6/x14SBLbt3wlJomBschqTE7/xcpw
gK7mnQ4sb8Vso5IIar55CN4e8Mr1ZYlHazjuqIHzxV1vBneuYU05sXuAAviuTxDR
nn1FD6rcZ3j1aELOfk5oY063DdO2w5bRsU4AZv1C37StIzBL2609JNCqakVaOkKg
gRT/HcbZ8FvS+7JnurTyjxNTzxNFcta2CHG69EHKZxN96IqF1OgGjCJogs10bzwg
qrik4D6pv5V3bSXvk4e6d5TZ+cQ1lVLj5G+zrzK/qNslp7Ids3yUnOfw3F/Zveay
t884h4TVamVYM0UC8pMWhCJf+WtJk84llvZJ33dKCUr8iaSgm9zWKOC5Wa5vWIkI
HK25RSBAA0rLAECl/+meu8uvJhF79dQoX5CUR1YYQKZm/VcIO+c0zLAYJB0C4e83
XHbTelvQ3Yp2xMCzeHk1HySB3wC7lCJldPNIdhQyGTf/qUleByEkjW9eTpRwBl7K
iV527tgMBEIs0SrJIEI5iVQ5iogrDQTGsZonwTGvjYfot2vd6uqwypSXRuV0YxDc
2/GlI2pLnopPgse4ygE7uUmjC6wNQlOdqa7UYW+JcjtFZ8ouJVHcZV6ORzl/p6Sx
22U+TBo5yaUd9r4FmuMr8I7DdcmhCJXYghsmtqwdu0ICDCOfAITjQ6lywx4cZ7PV
QQLsuNcG++lyPUKDuzTJj1iymeCWepgeKYEXV0sy0Ocl8JwLyaH4DDzg1IA8bUX+
UQCblOZkfpm9sWtVkJwl5sBFWCZ8W6CQHY/D4C7NE+UzfDTSP0PpDxGg1yTRlmCq
MXuMmmuIkxvb+H962QC7YeLS5Qksr+jkBAdDWnVKZepZoUik5HrPiUt5Gp/TEqje
ywfEdZbKuAZkLPNMqo7BsztVQpbmNA+gO+u0yNRqT7+mcZtykhll1AmQdQk5t6LD
KbaLsZZuA78S+bwMKncj5S9ZjheriOi1tkUIYF4Af7HcX4zWndITgO5LaqoHibhk
a68IRPnrYN3uyBcp/wlrfTskJc33GCsGriFbOrIe/ie1o+ACs4bsbORBSciivazi
dKXw2WS80C0KCy9jWZIpvoEu2GssEKMDE73akWp0C/yo2XLYipa1lRz8MZ0ZR/dx
QqdKW66Ksb0VyARHqWKrSGs1V9B/MXzWBsld9/yb+UfU4VfKbokHn3lTkpY94CAw
no1glTsoI1Czc39Qa9pBAVB9jy/otvaU9InsJ+n2HPOgB8HymIn7yscnW2SRi7Op
Br2Bu8DVAoIQ3x7nCb0WCxRPlIj5RDwFsDwdGoCyperF/sbEdJmt0Kja/ZmHycf+
6wFUeAKkf7kMvWWGKvvtbCFngj9DBfMj0gGkllYHQye+AoNqOZf6Xe57e7SatJL8
4/qNu+LXfGpWOAuW7411wK5Hhz2C1m4Jo+0/VhUb8zKQNoKf2MXgi2GbCHNCRhLw
rU9L7AoRMJSIA7pZN769Tb73mEccAR0KhjT0twAf9TOEYHbflDormbYcUtKwbDpm
iIOPshPKSuVMWgD8vW3u9qGOdMuIXe3gitYblO46V2e53DYasTlJHGJaE9EKXYMX
pKoLumB126GsljOrsqZC4fQyA4RrJrcG8CfEExwPI5Y/XlQw4PT/d5xhfUmQRRZE
Ro3/QcyW7R8v+ZihvQoKAvFIVU6/KUfwXmnAHl/GAZDUTvUSjp3yagzwl6iuDCtF
qc9NzvSuwsvFB5MwF/3hGAYzpqZkpoR0xvpSmmTXeV86nWkuOXb1Nj82hEwXfzkc
dFRtVWkr+RLGc0wmOniLn5Nv91gu5WaXG8FqdyYW1ty6vyehGSoLGGAMQQHy4OGl
gYjPjAaPeNvyGVq70m5gkr9Ru6VYdcdcAzT6EC26Pxj7xBftspHskAHk2vpw+JAK
1ESHUQfhQstYxu/vpu654SV94BOa443VQJ7j/fUKErgRlxhSeMrBqfwXsRLEaNyK
49Sh2lIPT4q4+4FrWYQ2sMUSc90+ViTXj6c2lz5qH7aElUMcSMBjbotQ7IGf4R6W
2uQKiiRyj4arkd21YdRkc/Ir+U2skiwU0qvWZrDTGXIeriETJ762wZs5UtB+EOj+
8V8bOqhuoh18fHxxGRVo30PgBDT/YJTpISnH6EhjEw4k4pMsEPAZGxVgUxfPdz0w
1XTfoMSytyoNlmlyXBoCZQcbdUVXMzYTrjAu0x4zCPm6s+324OfVHRTCGdnAgJi8
uxXDHvgrN/tqSywBSZ+RBkfEjgg2U5s0DLUSrUwBKrb9oWUJlWBxD0WP/NagboKN
sv1E8/MAYRZk2Dvxd8pslKUDUUno0ZgeH07TPPv551l9oKA//AudOrXuBhjXmN5E
VeYep/piENyGNf3txGyL9RhxykHk3RMnay4wLGFFuN0ThlgCm/dLQXHC9dkiFnka
p1Z2hf+HvD4J1hdrlmPRKzd+1RPa393Fq/mUjDLqSfFjva9XHEMGRsyhfVkXCN3S
U8rptCGqS4vzGxILBb39jPEChP40AYH3IUR6kkfz4H20juYGOjOhGhewREK18EPy
uc5/FNeeDHJPHoTDk160UOZq5uBd8qD8sor9McJ5sHDVo6r56a5jyKuAQHfz0WbX
mFzChMd3Z3krVwEKwiJLYOA3MA/5QsE+d6M7d9HBKTCbZrLOHi7l4kEPULHSEjMw
VQX2+anuchjsfkYC8UE+t+94ODqxZYGj1kGIWbnqmym9ic7HP0b6kTLlB7zwB30+
zcVdoEJaqKIH+qZPcAxFhFSKJyShWfiCHrvhZ1hVyruOR48YF1hlHch7jeKsIOWU
TQZIdGImfpLhoEr+qBeScJt3dJvspD+jvp4SOBf18ZIBaG3pXBMHsRgRqWSI3Pqi
rQkrV1v7NbPALmR31MmzmiVpVurtZ0Bn1Pwyarm0NXuzu4RLhgLLcndBPdPZxvdd
DBIK5+D9N0umhsaNCAPTTGsDSYilXdAB0dLojkyqIfuyO4QJIi/amxyeE16ylnLS
U17Pe5UJy9GPyC4FGKIgEtM8PNYyDg3ZQi+gXPXv4T7aHJIgVZIPvjxQVfABHtVd
WXj/yMU8QVBDi59AMomgc1271GSQLYGHnVhySy/g75LXMbvyRVE7e07UBdck6EUD
T3alJeeW2OsTL9Pwm13Qqou+EEvhdolBUaZ+jQaDRlTY64f0tImPYEdYuLqG+Q1n
/8bBXE7SmIAhc2/5n46pKjn9Z25G8Tj1l1HmbIsavpVCND9Hhee9ULyY14bQ+Vvg
p8EABg7TLgzPtEBizKu/tQCF/+ltrC4p8iOfIdRX2CRzvIl3hrv9gYfivZY3vKWv
mXjna7VSb/qSI+PVUCOOYZg6BE1cNgEVZY+tE1KHHhnwzPZwTMkjaBz6ukhBqKbj
FRD7FgDy460ibWjyn1jl+SDstiWIL5/gi/KUvsv55g73V6sz/A5mJ5A6fbF8Pqzu
JjU41WsVUQOHjBVfum/BmU1c8PRsmmw5b6x9/shSSx/VXCoH1QG6BW67Cc5ShjvU
PU/PsZ2VpiseTKCCcJhLQ4dWqDwq4MF8DL0CG0r3acdWv3VL8K/al2NKcZNCI+s7
pB/M8HTr2W8q5AFHmgsbCbZlXQs2UmuoK8s4GKtvk8OcnMNI7AGy/CFSbGNbfYbT
jEe+jlTHGakmLlkH4LEAMYhaSHWJ1/Zs3OS9pmgQDRuaZZuVKOMFf9GSZU5Bvqwi
0S6rmCsdDuxR/oyCrBLOTJo3IRm4Ct4vlgiLMdMMiZanst5hvlBOg27uS4jubHxz
E5j4/y/uqoHkpgVyeyYvFxq7cFqx/RjxzkA5tueMQzBu1n8atrXol+2GC1FPorLc
hU9h6Y/1F5h5g/8q14uPfI/41JigOQzFFM23Ei6C7meYRu6Jbqh9ilZNMqqzESyT
FxVTKkpYMyNFZh9fp4nNV/wek5ifPKggzUgTv0orMqpU6hzaZgzB1+/cdqmJNirP
bdvxQWHRk2xmQrCR8Og2vQgU1JnZhJrhXtAgyGQ/3CppOXbImXNPoeu6Td/Ah7nL
0UPwNb9Hdy3bKDr9Zkdhtn4BNHG7eQ9BjV5STD8qXNjM05BU+PDLzK62KqaP79wO
fZnvGfHKJTfs+lUZgYWVO43FKP+JH76z2Gi4585U3EXSR+pWJWMkd4HXVYfvH04k
5CR8PwDV3WVxBAhgA9bNxOR5Lh6irIblk0otZ+s9LTTxP7TFJqiyioqxb7MGcDY5
VbMyTY9hcLsnXGHfD1lcuJRrhijeRq+6UeexgzMOXVSjx539LXDNmsSt2l+MICY6
VFn0YV6zz2vKAN5gXUelRtenmZJ9Y3Jl9U0oBeN0J3ytAr2Y2HJdsK2LRIwyP2rd
Vh8zLtnSsFpnltsqQaLG1SC0lxYRtcxvO4LFtplZK1AiY/5pK1eziRewmKe0CdkX
KNlm7lOFtwm/lE3dSFroNXzUcGawcnBhDFypzjX4Q9dKWW88xZTui8VDjSZtIumo
S5qDOLxazYB7fBxSTpj+wQ==
`pragma protect end_protected
