// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:01 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VYvKXT7BGUBPQEsRTaayYNcwKtiloMVsS+B507C57TvDXlBcdFhm1Ezh4yvkmia/
SR7Zutki7GGM01N8SIzH5YQEc6gkIMpGF87oigqaV/M26eNHK5lBcmREpKgy3eoY
Po94gghpdObZuklsPdvH37x3djrR5sfHe1vrM8A3tHM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
siiZcHP4bw07tkdo3X3mZDInCQWOjnKKz8vExgwfvo7/yHfN6BHzt9p5YvKdJVA3
D0zySuMrmMix0aaak3o/Rypgj1QnyJGng9+LmIutl8Ilz8ufY1XY8Ptd46d7JfVb
kc9etxrVz9KZyAtVbMRNSYG6k1I8mPYQoYojkj5ByMqIe+pDnCrwEIXzMQfXivRm
lOg65BEw3XdFz7Zxj3uTWRVApPyiljemPKzVCdNOcDK6oA8Z1FkuKmYS3P42t613
8nHaoxuoISfPu9+kWAaX8JE7Rb1Z4iHf3rRsMGOdDkwEFALDuJN45ckXD9ZqCMk3
cVJohOhnMdDxI4PY2ZdVVJQ8BlflY235lwF1k6UDEB48wn89a9vpA7Y6ROLIRgJO
m5w+83MRs7LfYw8NvBkuDnh7OQ9e3ehpWiRhcXYPhPaJqfJllaXpnieIS86Ir+/o
5fgjPbQ6h+H9z14Aclb0CRtM2Mxl1mT8tzo9DhVL4kP//RLf2u7pxEOSoHWUPxCi
cVyA0jnbKIsrJ1P2IMHUFRRihHVzzK5FsAMnG6oLmEwm2GYszkO/HHUFF5uELA8s
KbNdIUehvADdp8z85RUmL5GxLhNmMDCtm7AEs9/JSeU0cveokf92CcbjSDmpK0kJ
Gw5MYtJlMHXHBxuBclT9kDPllIg2KzlM1JsgPTlr4J50H/9YJlRFWzYvOV3u4Wjd
DmJd62GAOK/HyXSqAElxr9Yjh/+Hjs5aWnTdMLtyvJxRuCZFwmKnK3WncHAtrh8u
/HgM3DP+rKU42r6nYYnvZr2UH8dLGQZfw2RTOV4OcN86QpmcOYOjCY1IMcC1D3Cs
ijOrFGsiLRXR8IeBFV1ZsW5o1GcsB5zoue4SAkWROTi6KoVW28XEGtFBNADJajGi
TGEcCA0Nt/6ZzH52BqCZq6bIjjlTW55mZMQyAkiwHuZQtoCvrZZSNY5RBWcZgVlb
suumAV6CRp7QJxxNpruSNYRAZeqdnKKOgx0H7HVGK/ztcZonDCZ6Bef1Zdwf8Fp6
QUTxCUHLP5iohW2z9MxP7zHo4fSja/y1N3EAqb8R+PVM8YbzPaAQnHbYIsU2I0LZ
r1XhnMFYAl6Nc6tbsoOQlV2DEIrRv1lJXWkEpvSGizbMcrMEqdh8fSj2Gf958UyM
VCvBSqnDSdE5Dy8hbgYgqFCXEYN96zbAsGukm4TfKyo4KLfi26kkLMQEPGnyoyVA
Jhv1R3MT0futGO4OlA1w8aUwXCKgrWpIPRDu8HkpfPKCHp+RTo7wIoV3/ITe4Hi/
pf60GqwbBrUH99MmI978DBUsHt3gnzDhYfvx4GBri1zf+lHHY66CNxTt/2hESk5l
ZV12XCjpAMdLut4q6hX9PTMkSG2lA4cUEvA0LJMq7j+5U8foxfCfcvPdxbkjh0T1
OC7rTzjx4zWCs/l6SBJTWfjAhJ1G9Q7ypTNu/bI3LxmYkMrEJXKGpQlh1uCFaODo
mN7BodZ6WFNJRCC2GcsUoM1ZxdmpeHpvr42JahWrYe+G4WxxRx5+JI/EX1qXuE3i
LhtF+qwXAJEl/O0+FPfxy41YVhtltaL9W98MaXCVLTQxVkl4u2FSQsBHUfckvuXT
h5a9gj7WyAVtqD8fWReXsgs3fN4iTsgunj86AF0isVRlWN3b9eKnp/4/HDoSYq53
HKB+0aEZd/NKoKlEuQsI1zckDcDrEzR6d/v1fcjaqLabzrlkYKgtQeAe/3EVnrYe
uk6mm664Ule93w+dZerpmngE8u5+DeL8DCOMgteKRV1hE0HK0aO+eXQ+zQalcuFr
a0GsRmc3SjN9HdN6z1Bwopag6UXCA+836l4rm7hgXWUaLG015SEu1pBumnujdsZD
DryTD6lRegavUtW7MPkUvg74ZCEbEDlfimcsDnBMDzs2nEEIZoBamfqfwoLHUrZ+
KwZQiiYf+xKObjeQZFc014kySnLq7d8zaeA8FfmMzNZ973fFT4PrYjQM8cSBXsmN
H9iIcAdfG7RMge3RJp6dbH2Udm4aNP+L1XQ+Rj9hG9JeaNFcvJHi24wyJpkmVCYS
zPk2bXIBasuSZni+kJTpS5YzpA6JHQUMzzXe5GckZ/QfMnKMLMlvjESkov9qguVO
wpNYOzd00x7YfHHz5Xon3V/LwxESA4AL+Jo9b1inQDXGiVdYCegVHMgLlP1s+v2T
+dw9VUIOeu+YoIocFnyKt8PfjHeUWXVFlLuzjcYIn+qbKEa7/kEGuzfkQqUvQtxH
pVNN2Mf7ZFp69rwkyNUCN9bfNaYhwyeG+xeqQXnD2cd0Pt8BjkjX93MtmLQ4JFyG
5BWXBPg4pcdd0FciQjhY9r9+dybEZtRDn2sBULfC+FL9uz6xWUjGpQvxk7Pi+rjD
BkglClDmfOYNvHVzw555cxrZFLim6UPNORwPZ/ksH0eZ5SwXiDMLDVGkgzCFLa9v
64yh8X6F0HD9OK6fry7YMnhKTYxf//nLuVDJqbyNDJ1RsEUVyPybNxh9S9kSKZMM
ylaX6IOJghM6PfRY9frrTyIkZnURMWTK5/ESBqaw44ks54F33ZVtnv2iaQiUDUOS
jYc+7ARL1+dfQEZju49aJ5hycQ4ZY7OShAaP1S9BfOY0w5FvxwGCTP3jZhDkOVJn
EBeo6gGO394WHwJ5gn32kTxTNoirOC4UzQZ8ZixMKh5kIuRLZW6f32XBDHr2yy18
Nn9rS1YBdXlRu5eStcIlhGPlN9Y9HG0wgyQflSU+qjRoJKxAJWeocybc2Ql2uRtQ
/J8TOAReLsfhk72Xa8LEHGgWCBscF3mgGvk6JsdFwz+eiM2jCXpO/82rtEc8/Vau
TEjGgal3Tf5Xhm7qmUxlrB5Rrv5tW7fTPL8AhOZDw60Zw+b5RiCvXxIZkN/kcXXH
9bS1CKjE4hsSRnKNIsRnNZ1xivtXZVLcxYy5M5dVpuAJflJWNAdClBFW780CovCh
a/zbiB+OVv1cSDOUFzaERlvEVgfZUTV0PDfsHAlL0X0o1sGmtHDrq6T2tSCYfaoL
c8a6XKKUKFpCRxm4Hil2CNo5Xn3vTsgyvu+hNwENHO8GuixP9IjNV6lBkypGjbtL
zo9ku9JcDbLHOKmEt/40OyYaAwAIaO7IT92LrH9vb/9N/H0CTO++QeWiZJ+HCrq0
l/0DFdZEz14aCcyU0YOUf3GEuZwxmXj+4schLCZg6z+imE4kXtfCaLi9MqxVzoQd
BFMS25/ixajOGYqbjw/C3FJcbl39JyRpIjVk+UBODh3TZ+UJ79BKwCgqZ623i/pG
5whWmRpX2b2wOsRSZvS/ny9rhg8uiSCZe2WnF7M0PvVrPwg+5piYrJUoIPwOYLCU
GiDhaxuKxp8sCTmSh1s5WMVINWFFZRJgSUfT6m2Suvi6oNj5byNfHEHX7V9b81DQ
1nHJjq4MLuQtaZaoBiSWQH28SpqBj7ZU2QZrRyQKHP43nFjY06D7meAPAkoP/EBp
EsDdI6bLFiJ4lT4uPe4J0aVmBXFZdchu52QKh9cO5fgHI1/iffIKxeemBFEgg87U
wtYRUF5vj69PXar96CMOaNnbBTqUs55JtMgaO64HiAiFv3asveoOA73TYUT+TF1Q
5DKB7as/jf/K9esInXHyUVmim3q9TAae7yQih3uA1qvgu0qjxebAR+imUuBihTb2
ZsGcihw2nzh75zd06lgsRTENDwzT4xTKApFyn2Oy6j+PbzFxuHTnzOplB3HFoqE9
YoURESRVQawE23Rfa4OU21TCV51uOdS0aoNbKarMuY+ftQ4sITBZB+7rfST3/qg6
1RL/eVYLBKELTorNR3yTZMHeHtc7ouUm/RCZSlSO5nqiRHTdUer7WQMoNadV7P9i
FjJcRiJhWgl7l+eD9hLyB3TC/fPz2gLzChCuvKcFJ9vLf2eLiAfd5dVxFgYohxuH
8kXzj4w7Nx/wYRmqtbFXFrrkIrJsCyWYArWojYEi4e6bjAx0GsK1aE8SsuGcGasa
sUPrMaNW7DDuv0sM3TepV//uVMLFcondH6TtEJkJBHxePs/2b5EjBZg2u6Jqr98J
Okzz0ipe0OkUHQiIrpxzi94euOCc6uIlw7lc0CqmpAipXOu18L7RaNekGZBpTavl
8QdXgiFZl71IoQDuffgnUXS+lhoZ+qectBFwB3ViclVqe2NEArumw3at/LvkOkCa
MqoIqvwib4hFoQRJSvMB8j6HoW3kUd1tXaDSKdYo9NvnZc0wBm4tETNkbIWkwIv6
MpTPUd7w5+tI0wjT3wX2xOtkmHB08EzV96OLTyjaonWP0zoVwiHkRvDdkcmvm3Z4
iD9JEmRvmwKejk9MC2tc1McEDd2X5btUFc+D1wCR1p9P0WQgHfDOU53FJ/GnakvO
53l226fWUwzKT6uiofEby9E7F/XMuHq7TpeXYBLRRaVCDQ7ylclEl73ffFvXo5dY
cVYQWWJ9aHreVu8LXe9vcaDhtFs8NZNawf2KDrgALKZyGKJA1Smtwllu3B5/aAEu
5AFo6p5AvG8tHYoPH3vsdbH9MUdIICXmLplswJGNrJ7+5pttAs0DyZ+kwlhuA1b5
wEevk+C09HkKzv4rcB1qVvvEvJhMSlDG0YLuhUrnCOHyOAS57JkBCFMs/ZHYbSDa
ITpNYUubX37alJlOmyrdTdpVIqQmY74pfE+kIVTiNLupZGL/E1Gkv/ko5VJJsOTz
ada6jJ2mbQ7O6gyLDxCAXVr9jzutO6DqkI6S26EBrMIBFQD4Zs8cuzNyoUbmcPUF
la7dulv5SvNmxDHVvcELVKuP6kyu9Uq4I0RCtb+yyGSIysamLNV0+qrDach6JOxF
avfoiRgTG8pe3JpeJqCGxXxGK6lu8+bZzfZ/mK/Va8oI6b5EtxaDXqL517KKWIjw
KOLxJLfMqG/FMcqMFRR43ar22efh2cR+k196HgkWKlQGxb3CO3quxRnr+ZjEN4ZO
tXUyBiPjo0yBYfD9D30vEXysHD/5JGQEInnugHnYP6xCNTS18+/ScqsOmQs26w2q
BI4OdFIfwxIHg5Bc70moVY5Fgn526O1KDFGS8CZckYOqwpf8wWX+bIKxMYZ/9zN2
D12IQv0C4ZA1FSqR5sbSkgE9NYeo6UOAjCrel6CyoPBfyOTTWvByzEgdTkOfUdBK
gaVRaJwy5YldipZ3CIJwfWjjXlq7O6SsAmxsxNYDSCgV1g4UV0hRiKH0D9SUlw2d
I1N8vYXFdDo39rcO61At5Lj4NuT4zqb/W1Uv5fuqrbsIzrL5ctueGGvkrxvn+O2A
FT037Ky+Zt/1vfDUrAsiztWl2VtZ4yzxM16LPKKQg/Qu5ZpjDQh4und69KZOJ6OS
rIb07N5ZkoNInPwyNY3etC1En3P1jrOkviYpWOoLdfTotHRcuyl9NcQ1KTJpePKW
gDT8OfkApF4Dy12f7grqun1qVgqHJc/UBXma+VhzwP4M+DZ/9FRtoMzwGoocShm4
R38ANXtOWpltOcXcYilboDXAS0sJLLWGx3W6JjtNccj00GZQmeLjZWBNsiYGDZwG
loTOgpyrCntPqUtkmPjHkeWRc284KwrcJ5oEHtEQmYitdkF8DA2k7xQDQFReclp0
AuYFm/Pg9STvBC7I50J1Qxsi0tkVdZ68lrJO9m30uBwWb3l5KF4AUEamNmcGSupp
KJbC4ISUlW0flbJBuFBHlaFU6kbnY/pxzdpu35Dc0ESKEtyHk7ac0iXHeTSZBXYc
q1V4J8Uqf0oZR7Rbcns8cJzcUBhovzb5p5jY6jNkJbqn5WI1ufTbFq5MH+QJR8FB
r9Jy3+E0uAkPC2vlBRQIbceHj7UqNMDI8aEyfsRKlrHp4CaLCt2fwS5Jezaq6lSR
Vgqtf5Aqku1M9GINfSkohEf/doNlw9U8nnWUJx8H3Kwpiyl/dxR3xGtpvRd5gYO6
rFLSOWs1ZYZUYutc7CStQIOny/DkV+ypR8bHmlkk0XR2MpxCsaxoahDzKMUtEfBa
d/5rSdNPE2ZR5QCj2Cm2Ztg7qoR5WWB1Qh+hwO9x/s/EatfkF/Z/zJWC2wVzP4Yb
ABexP7+DF4FAXpLKzl94XiLlWCHUIkevlzvc+2m4eb2O/AOGyKNqSH/uudKMJ1W0
r3uJieiPlsjv/0Fu8rEGFVaEVMpdfQ8f+k3AFryiZt8h9m4U9av3F/+TAYE1cVBF
BX0MbNzyZucFhL1IMU732ISReu/19B1AY/Eaq//kYOVd33XrVxDFZL3dqGufxPIi
5q0DXacMnWI+Bql0ed7Yu2ShZd91yM5hN1nhn+leC40Vgx+mN+aZRdTsBCjFaPxe
VmCntZBWs6X7u3artpkb0iNy1wnoX8CuIbiGaChWdhZPsSx0XZeh4D6LZBgxx/Qd
yz0al+/JGWB+juUFLxbRSFPK/I8JXE9XiBOSZ5HvU8jCzMX2Xrs/CfhxyHlQqPLP
O+6A0ZXaFWqkZRXCgYmgRVqy53q5L6am3QUha99vGU1W21IokLOK17fUkZ6XquCQ
rkGupJACeh8ZunjfKv2bWaIQC3djjf6zAJ3SMgR4XWSEKN6GyT3skOEv2iSgPFoS
1jMtwiTqEHp45hv6qj6CgPsigan1YsXftSgcwGm2LV8q266RRnZi6aWq3Skjam/T
0+rc+6IPTJaK25GCLotODw/AQAHcCgccQ3HIIk9LJub6TNyJQTfZ29uySC1tQDV0
UsFDkpC9vERMO3iwdncsjK/buzNXCxAB0RGpmhRAa9NLTFbUXxlR06GwDedjn7Dw
D2Nl7NCp4MyzLvulfkzs1FpK6HPp3onH+/FTntLz6Y0SZxf89P9s2A9xR3KW5VcI
YEahc4a6Nv9KTBRH9eNQhqBmDkdyf+2epYHn/vLIXX1cHVgvTh50f0NnLxgw1+Kd
lI40GWIZGM8jdYxQdSzZSonJaSWyFsNVX9pTK+HPEPjCLuJI+6YFc19QmsX5qn0M
65KuF2pU/QG7jcBdS0GXTRfpz/YSY/56oP4FZ8L6KmJeBQuaziQYPzSCJX8hFyaq
D4R/2ffxZDl8rthieydKxnVozSsNO4yZ9h7wdvQNz9ON3ddmUMKWM22EWh8U52KS
KEvVSawWNQelH3aRef3fAG9qP8YG8SBQCdtBd+MlGgaIPS0aBKKjog9tC6wplJBG
4JTCrmR3foZy//fGE9ytF9/MiGFYFVq242tgcIjF5LZ+jfcHzc7kDf4JfTkH8bxZ
cWB9RaWtLiv+EyFxV3P3BuuY2/MeGg5Xs9K+fZHqLlnCyb5EwGdEj0i8sVeCpCnu
w7pSKXQogsAiTjrJj8IW/IpM6gJ3U1Zl1QzjHY2F8Sxn03ypYgmvXKnkOiuEWoAB
MWequ1GjjVL4rmA65FDYgBHOkR+vGlGy+WP/ygEL9WY/3/lqxyi4agNMPwWzKnBd
EozcbcvbToA8fPjD++JN+09+nOHW/Sk9PyWVnOWCffjWan8P0eFesZMi5QKKK8tc
CZg/wLt9zQwIYvd5pcRUMCMP2a0S2LNPSKjDB1PsVYVeBK7WG2Bvsv3zCU0HhoSY
lCpm4UG7sMquycGd2BAV9zM3ynpV3oE2WflwQgZ6K00W3Mdy7xAOlyMS//cQirXk
070uruueQAezcjhw793R9tIDIXBXRsMtWEKH0CBajLK7ulB5LSzzCBaD4lKRE/Rf
s1zIhAd9uNzrZEwLMVtt2iEypFf7wtBZmnBERkEju8EemVkZJxgirGHhFpeZJvIS
KpZuJx7kZf3BgL8n0oKBrYz+N5hlssjhqK6lDQfOfMb3mXiUkdgd2geXcsGX1Mmi
sDOGC8Mi0yECtf97auyVKDYXXD2kQDyK69QMGqnSrHXVvjvhioYHTm10fkpUMQgi
yZ3ZBLZNJgZ+VSp04j7Mt6ExKTgvJeUjClZ4B3kFDeJdtAXNjl5nrPjTT1RhLPYP
VYo04dCXMN3aZsdmgWL1Wv87xPIDpiCNNficygCzrk5nXhp2+g9JkXeWjmePVQgd
qk7j3feaa+HT9vWcRzuboi5zM5ty/JJTJK56I2OCzqbtEUZlt7z9NodVKqrJJ9FR
Y+AETxFzje1BycVfzToIBWWZ0JimWGVf405ARUcuMKXXqW/VH93daJT9VwB6WWe6
kq90t1XLGklPjTD0c1mf9OXsemzha16/0m22IpUqokKzyKDuI4vHuWYb7QTHU6Wo
e/6iOf7uS/2CrVwssceU+gmVvMSIfHW47gjyAnh+UxFYai8bOYkMjkJC/94g1YNE
qob7Z1neOYHunyivgLSSGOWYig6JbqPOo8Nf5aG2NW4D9JeQLP2Nu1XsbD5b2BVz
GVidOWQYg6lY4GknUKTj/XPwhmT2NMsBEt9VeNu47J2mmprMYgmtRAgr5guwNBG5
sO6DeFYY0Zu7th1POgVv0q967lDrS2Lyl19TEqbSpI0V76KJWWGpN1HUgOrs8Phr
8DSylOyJTdSQjQUfiax8PRGZJYk6bT6Jvh+6bEIaIGrtBVSYQJm2YYQKGLd41KOo
AR8W2pSwDgN+VUXsxpVf8xum0Wu2XoSpXz4Maj7sZLIV/GMxFw4IU0WAuPKab4hu
ocy4+uWg4KPNKDxlKzEWQlpIaIW+zAoJg2udnvl22Y0C/xpb/lLL2xvcDzS9qShd
eoUTKU99DqzO7vq1RfCAuuv+Sa8+xqGsfNRriVdyjNCI8xeW7Xm1izQa3EtaK4tK
ffxsnhprff51EJJe3iYS+i5dAzKR9ypHwKSjXQE5g1q3ljj67cfsL0YYsPP+sL8D
fcTXw/FbC1il6wM+xTMJQp+f5e6OzGsfClvlBO0VH40PjeqD2F5qdNON6gyGG5bK
mXn/FE57/12m/GKAI9l1EX70yqbOPmkXCJbt9tQJtuf0q8JkVw9ElnjxX8836pVB
H/9VoZWWfRttvHUBaZKbz7QTxlZoJ3dl97xUkPMkebw5/TJt5RhOvIeob1yy1Pmu
nJXcXThBDESanfrufXQfSARNYTOCOoyWnVocIULgjYiipGpstvNrIU4WdwmUsTTz
TiDyr+W7aO2IzZHWDCEw0ukLvTBIMUnqYNSISVJGeLZMtkisCWlg0qKd4t+8R9X4
1XjEiw5p1j6uLWsKwKSCUQDqgVY2Tn9qKZVdB2oX5v/VcdgILqhNqSPl9swbfrHK
9kB0dH7HTGnXX7u0HU4lQBLNv25K1Ygn0eGNtjruKuY+g6yQpXZkuCQeBqKwXMUc
bxT1UuZjsHXJwZforpK3e8LewXgLWr3dbu5jbA351hcQ+1Vv8VnrnYfOMWQ6yURm
GUp122qkxp7bOckLCpq/fxg54u7Z02tv/aI4RbQFuY45FjC9Gq4rMe//fp31gdRa
+7vzi+yFRsJ0QN7lBAP2NkOpdjAJPcqnk3aQnKpCPL6knZ4cgYs3NaEk2CyDYY1T
Y6/z6yQK5j5xZxAnSwPlOGXi6Tm6TQnPXNTZkHHj1rvjDTVZ0H4H0pjEawo5sVjU
qaLWai0xbz0vGSR78qDEPt8oBlsHQtqNj07ANJ01EwlNoMa7Nt6rccc+13CxvcSS
bCy6FKMZ6Bfesxp5vavM0APrMyh03alaXVsKQw1R8gCtY4aaMPfvl7Ew5dybkLWs
TWNLk6nGx44im28aGmq+ZHYXhy2sb+Qbh4cPQFvzuN4mfGsfleMxm/s5qJAVEOmc
HBLiv03heRw6TunQ2gugZrT2Vl/iTtVd5Ig0mQmLPrUxek/is5u/4HWc0DtT+t0q
xuSdmcUuAsqv7yoZvJ2058dIjW4bPcx7ULqLeHkCPXcIswFf9j2p1PHwqaeTWutG
KIMyBMdWZTOCQv7usmQjU7MFea7qTbhnzfHgHgKwRO7hn2LcFJFQCy2e3cME6HG4
RiwUPBkQZ6mQAt/YF0L/SRCaIqPGUbjomXWYtVJqD7rz+Z/Wfrm7eQtUBxFaz1wF
IGj0A+ior9Ia2p93s7Dzbw+vqOJBGqnI2NKTqsr3P7LZgEO7yirCChJNeesn5ru7
n9AotNhKh0f0G+39jbhZUhI1mlSLXq7Mx8V2I/bM7ABiUrPqVoQevFBwvH4j85mT
SQqOAVh9ZuC821wJK8S+3MZFZW/HUxtQW+RVdFUGMfTnksbNak9WnxHuI+NJuISq
TCZhcN+4y0Zh15TWxAcjdyt4fyeVGmLEH5cEYVtmoJM=
`pragma protect end_protected
