// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:56 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tZVkgQw6rVtmPpmMS9OnMkVo9VEsH1crpMikLOIDSh8MJWv4R+Y8h0F25Jx873Pj
L9i/dknJRtgVoefGJ2OcU1q5P1en9hULZMLdKKGk62435MOVNlZhReNwAWsS5c6J
ChTbtGzryTDup8JHNcsysQ+XmbnVmIITbKOiDtzzpME=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
fThmatLOGTjiq2+rAP99zm1GZ4Gn5HgaWx4Pioo5QaW5soRj0BOj81fhTnI9sy+m
5uSMFhte0s8Aaj7SS6+SBErLQ+R7kN45Qx6aJZm8NseTOsDC6sA6EH3LplXQMz1i
IIObVrA41Rvs9stt7OFelBwtY8qSbCEP/VX/F4Q4Q8u8VGWkvK/5T+CSP+XvG5n0
8wfsfCkM7R+FNDsH6PBa0MZZWuL9bX0EC3cmp0QXCQYArs9auwkT+0ITOA0oiFXl
FeI/mAKOi2cyeW9YKQXN3VRxisbBUzyzHKMxCc69kPrmGH+zUiLfReVo04gSapUI
gdO0gGI8qsZJhIDQyptk5zUN3Jak5Qnngm4jfEUAEwCHVjUAcQH51Ccx2I+Oi9dZ
WqNo5CwVWPGZry1zgK8nvuPTubYqdYFiQ6CSvOrMLvqH0r9QaISDHTdnpH/7m+HI
1KK/tbmD5ufiCWT/dYlPRzZE9UNuBlGFrohTbfffAv7DMLgTr8EQu8VhQ2y/i9gq
auYpJnWOumJKYo2W8Fv7mLS3KDrqG7yvKT2igj2QS0CJ/ko3ulTQnDVH8bvu9n/1
iZdIB59SuC00zcSWioMytGXaxbshHnpvDkP+QuLyDx5KLP3vdN+U1JszMWuCrpHT
tpFcs7rNbrG2Fx0VdSqShopAQjwvDZc8+SV9LXwwqqwq0xGCDCDtzw/q8d+a2xlS
8qvmVLoCYpLc79fXY/8Hx4FV9PdjI5wzM4c5OhAzuXl67j0AwGEfIx2tnIU+/Orm
f83KrGE138Oz2MS0xRIuwsP8xCuZoAb99K952WIQ+yJBo8q0hUJXiJtowXss5eWU
BVESVCUmNsOR09AjC7oa+sAITcQCHzmxglyokEYnNwehe64DOWZRJxIuEimUxLmx
cBPcAJ/7Q+TsIqwA5/wa49xumk3Q/hjgD+Db9tLpIUE3rbHM88LVtufUOJNzKsuA
GVP2MJBkgQeajWDWO8UFAQ+ae4Ve8m73B7zQug8g6Pd/1TYHVGVmUFHLdTfAK6st
dlxiF0IZIwnArWXeGlFza72bLAh+/UgZJ470NTIzJ7PcZCfl7V7LasLSoL2l8uds
0RtfL5gQr0YykmZv5BSz0bP3Cb27fFzbLaEhrBC4J0Is37KExb+u3tFBrcKwI4p3
2/NvL4Fnjehz3Qaskb7R1x2TdixyHGkOfjFSrsYwl5gK9UdArk9wegH9K+Y/TU04
C6tOV/zQ5C19FrhcIxIgV+IMovMNOYFDuaW1hQXplJiXtRZli5gm1RfT5RvEEfJv
lpXF3GXMc3R7zWNKH9dMcgRhi3FL4J4mA8QrLVwPZ1YvhgUgEMyKDiw5w/QmxA5N
lkbpouMrtt+xDAr03d9OBc3CQ2IDdgcpUHbnp2AEhbWqZOOGmTMCZtT7QUdfsbkU
j2m2uGx5887d5Ac2dcrIaPOa2TmsTyXzM3iFHmaizyj54SMWtig3XhYmcal/01Ia
7cyTk4nghQ5tYC0QTbwqujB6SxFNwpu9jOPA6rzlNlpuybvdZ6wCCeUTqHSNeWX1
GnIDHMGyNQ2iT9eyvJ35dmCslWx7819/VmUJsA73Uev/DF7Ac8xdbqzvT0BCMtfO
LTSz1Y3LSyHaF36ALC9Di82ARuYuQeF2AW+BkJ35ZONC/JCna1qA7CcOUJ1h5Z3/
zWv+dRBQzJTjbCDprT3I1F5nVBAg041x3peBOAngFH0rRqFV/6F0LorosoKAO7FE
2jJkxSm3IdIZAJe9oig9ajKh1jR1t21Kp/7rDQjwgykvpIiKrwF2CZFE5S0VvUtC
d5w76eEJcwJlScGmGff3TG3JcM1xbO251WfgqXnGL4EmeiMffo1y3mtwWn3TXBCV
rds3f9nujITYLucqLXpB/A7cl37egBvYpO7BrdI2YjxriDlEOBxE5UpBkSYbllBt
1rQJH+ZOZ0d9Vn1RBqHg/+ftWIAjwlZO6DzuidFg/bS7zIkc8XdED7+9mZ1M6e3f
uML+b9PNFHcDJOxIRHgzHboHGJCqRYDTImUwKFTxDbFD40VZuDToxyUjRBv0Lfh6
mRG1MOcScwWuQryr70C7HhpNe+rw9xiiNPyl+TWLxWQSGdjgE06TxhmQTh6O3z2P
wDK4+IkS9VHn383Zp7zzRKqR1YJUGAvRBJSmiWe7IOAUDrqIvEOHQhW66j/m7OHt
WX4aS8xjsGDvOQ7VSv/4pLPfPUM2YjQOvR+1ADTPHVts6ApAr6875BFA+Xs3yiCm
EX0g1UBgaqhxcF+pPVp8/bCSFU4iIIz16z+5+5iu51wzClsSFTOAeb5AdSvqd6d8
/jysCeLlrMV3O4xOl2HcBZiVpopdhi4feaQY6WSO4A8HKCfwQnSnSpNlAKENib+o
Kf/L7FhwL7UMWbXKgVyE3yc9gvLZ08fgG/M/qt1sC5Kt4GEujsRKyhovtat4wskX
XyqKhItYJmPaIMQOv+RYcu43PQI0OrrKNBpF/AIby7y+6uZUJ+hnglyCXRnh4oBi
3tSC7NnBRS12k9SPu8mSLp1bRjxW7Nenthex6Qp0a/ISg67tCkURApF4Fvib15FR
m65pm4Moe+2tQflm4fRjJGqF9N0eZ90oUSQjX8PH3LtuiPuIRNaEdJnAoWw+bpjg
sQ9Esm22IHEGhAtMc2YJ78esaEQ790Sy5arm9ykQH/Gc/dxW37K6IB24SajwjMkW
8FRhS2gmAE6LmCp0ghRvHrimqxMvJ6rEHhkGyN346xxHu6430c/1JhqepcRRwkx5
wq1quLzwi9Zd+tnrTruW69etYDrrMXPCrCDtbevoUOtD4pWOBUyfCBfQBAu0EMZI
MwwyIviBvYRhuhhwLkWGuRpXe4XYJk5Irva3/SoQX7EPm3vTpykkN4wq7oy8ZnR4
+ZY87BFAwXcVUFl4zbvttRQFoAfiyJPKO79KEz0g2BW9uSaPIuz0ge/Tud+CtyZp
+KULDtgJ7xK7CToevqFNUZez3AfjruvacHIedZJPmMXPQmlduuJIIZFS6MyOt5Jn
R4ZBI8LtbcCoPRB6sM4ddWkC6M5nbttJkAyDWQDOcuRErNEzf/Z1ZOMrr4cweD+9
Eyuc+NzZLGN/THPHrs+eNCS/lL/YYlR5rDC2x89atUulD6A35QsHatjvn8LYOH32
ECOBSHKTFxLXXNgFxOuxCdhDji62vDFkHxIGDE+EcO7UQRhAFWomez3WUbZcqw+w
W417usae9ps3LKGad2ByjKMe/RZQhXPGRYB55+hpg5qWc9rVqXCkfLJUyskNQLDw
jhqENo7OHU7GDkfrKOOR12U20poYDcnC+DKDZGGyAQeMs5SaFKcllLNLfJ7X65/g
FPrqdVQMyo2j8Ki5TJWaJvVZjexmcMu0lLEvKdm6NYFAPpr7oTPUP+RkJtpkkd27
O5kJvMriTbKuc6bNPgURSsQrxjtMxxPr+vu/3/iYKiaCo6Ri8QymM3hA5Oy62gJ+
z7C2K5xw5jbJU5QCR2A4TmwyzS4J2CP/skV0GpAdQDR6seyQOO5F15DDrlrnihLO
yHR+46/l5YoV2X7pZw/rOcTyiWP7obEbUSA5+EGRjNy1DfT+t3Kc2kDVYbOZREqA
kExu4Upr3pgfxL1SsxcMzBgPXYim0o/wrwQczTs7mghqBPVR1G5M6ZA5Z9PZJTc3
eR4RlqKnDB6aep64QmvrcIFvelzwYflAZ6poGbq2DVu7dI939TvbSEH9X8JNNqRf
M7UEyi0qzUOJkcZwTJ0pm0HIKKoFMY2roLEKHqpEbN9bwzqH0bb5e6gtLazLQUaz
XDS1OWGJ6KNLNea81s1n7FKCLuYVDGxiS8EW0g+H8C0fIqvhaGPVr1gmvLXFzUJw
sNH0uvh55N/IuZKEU6M67ALz8sLThJsS14KTlTva5kx53M4/NrPFXTJvayxqju6P
5BRfyVQX/MLJVl5d9rTEPUTC/XRy1UXHwKGHMgkFILT50hBMexm908Cla61nCZkR
zSGf4qdnOsi+zgGPEi0CPuCH+ujQtTpfOj8//dBEdGgNn8X7Qb+2OtAKhWcnNQOk
KlfeE11t+cq2xvfktrnmkpLomGMOVljgHdOFJdIupSwDMLeEzGSOO8k3BlTjdEBx
syGsgzHJvmuFtBXMHiS5CQt4hICgp0fmHB66DGtnrHKz19GyXVsBu6Kr77IPSVN+
b59HfSxboY4+3d/7rke9ehyqFfPkqFXrUFWSUzBUDEF/edcEqPwuvUlZUM5YKeXq
RYaOdivdptLeCX5svYIz3N/R9LbRvFhm/fKFwrkZzVgfEqj2QoGIlLX0DA72x2lu
6HgoAcrGPBbFJ63uIGgJODnBH4qdzgE+u8k/oHWmjEI1PB+cZciNMGSgJ6WmFXtb
h1I2wc5B3QzpslwwyQWUd0tuRn7TIIbYPKW5+oWZXe4FT3WKCl6qlleBQhJjW+EF
D9MJqqcAJvrnDn/LoqnZLFWJ1Q39Du1MebHbEFffOB+0/RaWe2JLxr51mX2uZGVE
9kiJZ3sIoFAGMtCIhfUZSn4fhD1KBEHbgECDgLKOcadGUjoaILtN6sBb51bG/eLw
B5yX9quzGypGQlA88zoJP+DWjIBwSKkt1SdsjlRBg7+/JDcchREnFAf5pC2NEPqA
vqaHDK2EZT4Durs+etp5ydiXBwzEKd/a1QLtXKpRhmQSCROGXtnUD/+hVI/f5n0u
D+rU/D6RgR8KK0axTZWJa4TJHI1IL+uzEaMpYwN1KN3KZQFeyrQhrfRllenuxLMn
YsGVoVQC9PYgKQLYDrZyf8vo+NXrPpj5sn7MC67ljEXVkzMHOwA0TxjYxOmpFyhH
SeWYEjzZWnn/pM4Q/DG3NUxLMmnoPhSyJAEZqpB5B87pjFkGViL/cwNCt++0VMg5
DAM72oT5TqxC8NFnWM8moIxysfqSj0au3aoA7BdVecHdTXGRRwX725pgjAmcXufV
+h8RSecEqDvhHPnd+0bW9sNChDtDPR10BvHzfaPc8ESjTyCDO62bDk/zZ2emU5Q5
XMJKAYXtO20uX2i1uHenJC3RPDTes2pPSB0EoW5lHMGHAyumDpBSMFtbzyi1WgQ6
RFuihy+93+eFxm7RqaB9j1mTAzEYivgzqkcF/bUCoaqTJzxlCOVFauljQczTgGo/
tFoaCkkwg8Ej/8mwwsTQ7Bwf//fcUs3eDJtXRHKoajYLzdosHKwZYhevyGMRUblt
ynHAC8Xp7R/OIjaJzS8d6pxVra6XizMut3RrJbuQJCnTevOTUZ8Il0x9Zs6q7Wn4
3ULN8BXAfXV6E++Jr7MXipzVVge2ISk+vUp9OzcScH4Vek3XqTgG7KBBeUXt+m1Z
A6EVBT1k1vrvEGAbTjQlNS8FgbYwP1DRYF0MmHg6V3Ugp44/u09OiU94VjZUZmxk
OyviVR/eRjRmRqsHokq40VZpLFLCazTLeDSDr72bcaYEMV8JQUtWntkE+slS6PPW
0vCdc4ADOI71Z73hbDJcWRSzGDQ13MMRnJe6l4JX4jfw8dM0EwZUZ/R4FP3K29Gv
8WKLIendUtOcCy+s7f35zVTQX++ZovC3fdXy0xDzEiZ8gHQZG9pLWYcw4/fmV5t2
B/GLZitTRBqXxnY/03zlWyMBVX/xtR6oOnUVITRGCKgsyksRoNo5usq0g+BkOQk4
5aQ3v1ce8cSIvKhwuB3yNCGtCfsYQ2YgEoMH9qxIklK+tpw9F8S2k25kX1hJR0RF
KTl0rAnB0iFEO3YdN8JvgBFpDD2+Y2mi3Dx6vvC3vH3T+POyUNBaYXVIbQtpBSBn
9ujMNbbF7CwbKNGiGMko8snOurjJL8glUa/BBut7fmdR3clXxGHqLUObF11XCFej
OVRKLi1LatGdkIPK+HLWIP/NGpEOdlcj6vuRjVXh67KczVrcWltZYt4rsk0hB6tD
cpg99QkX5Ji3iuBzSDe3rx0qk03KtUmktAGBUVUkSemOZSQUsxYAwT+SwU2LDiso
FAQgXJ5r2afVIEzHI0UVPk7+Rdrz9kMk6LpdrFnWTuljBL/RzGPmj9gjn2TgIzJn
annHn8wFGHVg1AUnUe53YoebZe9lJJ6mrjiXdqRV3YHA4nXZorgePJmAjGSSDnLW
lnz9dE/TYdwl6Bw1JMhAABwSb9gg0a9M/EuiX+qmM3zTJfPD/yb/Qe6+5rCqfyVn
Rm7nHvbPdtzY+5mZQZF0yfWYaDsR5EWzmT9EU82hOnbd4Q61R+g0WMNGePz5wRsT
xlHz45PeU9zR/cAWXKiafoN1mAL1Rxp+yQUhVOA2Nc6J4X3ADUIGjcJ7sg4kUTzr
vv8TSARH6lvxCLTV/S9D3dRyZlRp0P4COKirtE/TZkT+j41gsMWtJEYLMTsxQF1m
zFcAP/1tUtu544khQjv+yP74BIbAhtKxIfyVtzSsj+U3P8PmUh52oYYv3ZlgaebV
hDKI+2IDw2YlAtWWF03YaYgnQEhu5wb6lqRi9vocC4NxmJLyKT4zaLxXcBmUj2Yd
Dff/qw9MpG9ybuIa7lkXRK3o/z20XPIv8QBUc8W3KECNEIimIaYcrOH6InmxwZJF
b/8OzYvK2ksx//AF5wrlq0Gz4gFvpNT3V9th5k4k6qUtlgjM7AToVbLJpIgqpIxV
POJwC43YJsQtNaLtpkcvhSP6d/ccfAtkcffj9UehYDg9fJn0QUje7Y7q+5NN96QR
cw1IC2ZV/t5lxG2EnBelbiLHgFm5BxIGbKQAXCE3zzgJ0YLax6IC8Esuj6Xqsg/6
htC2eFbelQMuFSAV+ocNuHAis4Dbv3vVud4iY3Yg2RX4acqF2xF2pDtI6IfkpyzV
DFzji0OxwxaoQiIbrc8FX1kRdqkJLvw0UH4VUfErvyDZFF8hlYIOeJOsoRHUrSFC
QZM5UyEcXzmJeMjOrI90SRkfFE1sMNgmpHzA5e9d3UGIjFn2tVupbmnbwTlNBgMu
EULIyDU5pYax6L9Se51MUqIwV7EfXfCtD7MleXH/SA1ycsafroGt8KymM+9HOele
6cd3WecLMYCXB6jtS0wGn80YAOxWvlRGN8AwyxYuybHpuLpHIv4KV4vENw9LLNGI
8fR5/cIi91zoUq7vyPtlC8vp2/uHVo6KbPG8YE8sRYrYLT+JPrnvwEp/lAFIwTyC
jfEWdUmKNCyMt2QOb/BXnqrNSZxbdSoJ6SIsZlKVnVmOshcN+5B7N3cq0Db2axZG
16pXyfJELgDZO2FizoNj8cd4fBjMJfdTnIMDxtKuvZIxPfDnxfvncq9PVUCKCBOY
Ako8pjvfmZW4gJTDpkT4IH4NExIJLrAYDISSwecya7UnAwQBFl9z4ChodapycxBK
ys8EkAORZYPios/kxHGU8JE4RR7eTq2Ac6X2fdS5xKof1qJ/GGjDkJhDdertqm3m
K83MMsRz+Zu/kCFPBGvXhxS+3zih0ucjd6zregXY4WZvDyLwtss6VkHK1uc/SWA6
XaH+Fk2cYhyU6yqrtRJnclw/YGkm1hURFridAMx0IX8miSdIDt2kpJmAe0FVckPU
lLUavkR1fgswAVwp8wAHM7ivyh5Tx33FzF7uZQAyY+VyqRoWAEx0aAngv+8fJ6gb
AsY8bAeOOlaFACgcxCOnEyX9sbYQy94Q3+5CS29CEp/LbPCY4ESPT7PJ9dDxgpPB
fieqGrrfmQVqbAjPjMayD48JXa6QabT6epj9nmUVFRJEWgXdTYz3Cs4UcoGo8Io4
UXsuGKJZ/fQMaiqi7biYirYCbPIIn1m79PABLQxj/k66QxSw/FJ0CXVNK9SCXQd3
QzleDiiaaHbVu1l32DvpSpPg93xzEYT+XuiVSQEsz7eMEwkT26RLzG5EdOCrGo9z
ndDzjwgf2Joa6k59/2J76j6M/0TNbbTGi4lU5zbvU/hxg+pmM0mB1mXG2VlPd0cF
yM54qJQk8Qxpmo2nQKiz5/zF4IUc8rmw5Uz2l2rqB2zmmnoJ0BPifLq+nGyt+d8j
Wr8M6PZe7/Xa4G0HkdWJIfK0b8Sg4jVMZAt5oaR6qIkVqkzOo2zKEkh5MZ7NC/gp
46euix/R0DmxmFA5MOlj9RmAhE/kun2A8EfRXBZcpTJEaxicxiSAjj7ZxetfReb3
jjM8IMJP6dZoHz2v0/jM4ri66oR560QohwAI5ConS1bSuA9myF7RjZ13Qx7/L1EU
gOl+cNhfjIaXJXRwSvyU9q7ZoUB4I5R8wHduVaEghkyXxjT11V8Mx1znmxjajoyU
o49zcdW/+hrw630jmMg0wwxQfSpmnXU9+IyaYlN4HJApmgqOZrdchn66iTDZuKlG
YLiBSwTzeq1h1AphZ/h5mCBplsB8H6YkVjj+Xj69OgFPytnY0U2Iaxk0Bt1MwS5A
y1yG/f0OOcd8v3421E6kPzkPAyQDQktfFkKg4F+MjLyMBABWh/ricPU88n155UG1
7HnqfsdJr0YpEm5LGwox8RJo7GX5305WsK/ZtenHYgucc/2O7HGXr4Yec6R18i/I
zCp/kvOdq6MTV8rCX+GdINP1HwOU/Yh7nrFh565rnwmNb314ISWMz1noJpKSuyDQ
wXpzDWXdiO3NA4OuT4ff+LkPxWOBLC4l7ighrAyS/WkGjLMBQTri+S5Vepl+SqEH
sL9qislBY++OYOg/x84nosVJSGjqqFBkSpRLnoTsa6j5U1BjU7/5ovmDpZKZY2Hi
9wLGxHRdB2c3lbgqBjc+MENjgHUbAMR41xWktMBtDWNFPlzPzjmDWdBCdK1YEKg9
qs9/g2MhjMTxVjGWeMARHTBmIeDReZiyUXurbKmLKTkaljpB8+VT86N9nvDyp0T4
Iq27GXsuWPmbrrWljPTg4IdNFKlsfdA6sAv/GxqKjtl+XV3451E3L1BwlmBH6UZO
VAqubU8BJFeIYy/WVEiUNK7GagdQRw8Zpuzqe5nZCkOxNPcvuqRTeGTyF91Yyhsm
vmOL9xjZ0sl5RAnEXLz7R6AFVmhJ7ScqLIfi1+O+Ny5TcaGeO0JzU7EO1qlrlfyu
j7iaNHKYQxF3lC+7j0Ib68XqZqzVIWovctd1TwuycdY29oRoA3NPnRbRKhLMzCHt
XdkwYIqJiJRlN793mA+7oEfut805T1dVW/c1NgTeBQOat1ZM1PtrPp3gPWZvwgp2
N6tpQDRj5hcVQ4uHOff43xN260qnVSz15pJYN2Rs5XztY1jkpVi6iv39tODFFhlz
HGCXVXjGbgyO1EHd/cF7nE8bSPQYQo0ibz8/9EPuwbqJJXu/gQgJjt2OwzpZ7xgY
eQ7bqyOahmw+NkAYOOhwtevu6HrkwID+4Ymsu7MNMRNxQe23Ddx9K8NedF+JYLqr
QcI0ExP+PgDbUJ9ZV3UEy2IbnYC+wsU4EZMZ6GV4W7ivfAiTP0Y3FxsHy+c36xr6
Qtdh89dxgGYZFOx1E7ogwAE1OmaKLXhkpZVECHFDV92mOqaFLP2KAyAz0OKAO2u8
DmhU4FBSO5VKha5vvgdvNktDwApOeVZer775EQ3bKfEhR1E4eDzd+7KvPCvvaMtO
7yteGGzP+oXhTyXir5XIZq61rhYNsOGtUBKHSVzxoxutq3fY6gXtjwLJ3BZdn98V
sep82i/lv+rHqRNcxF9OpHxSJVR4psJoVnfKxIBSSuHq6oNO1kTMA5HvzABM7XPr
bwOgFPALx60rQ8Jbk8xuBOnRiXjTd8pYl7EOREa+F5bQBY5ZPozSwRzMbPu9mrrv
hs7qMg/Ps9m5ZWdYGsvCewjBEiLNhN3C2KonPxnSBDcvjWkbwDUYP12cabEFEY6M
Sdc1MUnVK5mWCzmMsBTxnljSHOyNdCoEFxumTimoy/QwI0KPH+Bxjl2WhQ1LSvXP
wRYdurrvdx7fxrtWytAg6/22cCNi29YWuDGH34Gezd2JGwXdZWukgjy5gPQEPSgn
uJc+x0NUB12hkp7DyxMq7nOUbf6IqmlV6URdvMmiRg7mlB7UmbnojrT9Z/ZVXHzd
TkZhPFvRTv8KsT3Mt/AmMDGKG/ptDxdY4PucG/W2U3XA94Ew2j1hFfsG2YJ+aFfn
WpPpf/f3isCIBhWCS5KR8biOtodlCrSlAxZekNuNKuBPtIcMWdhkg3CG2YP5WW1Z
OIooj1jzJQh4FS0sRxq1XE2/ac/X7rsrRdrPzXSmqI6S6X+z21R/IgRgUTRBFcFB
B2CX6A4NqJ+J1j87mECtwRbZvt3bG5/QysMKnTHnKMhJZqbJ1yjvSaL3VeJvv7rU
6rkfozMMpkmhibWPCGdC4R45NdWHUSjJTPwTyeEyb0bQsli7Xom98F806iBgOYFH
HgxUkfvduv30P+0fpxnw4hJAuMKbsd8W8/dHmrmqktYjLH2IKf1bpm1lLzXifUh0
C2vxKGFk9qi2VtOLeK00mR0Ap23jinzQ0BGmV/vZ8SM6NpFT9dUqHjQexfDxpN6h
GW8ElWNT7SlNRKWBm6kUgfxlXeBecXTp5oUdu+LrKXyKCg3zxvddDVIEkLg0RCXm
QLJMLFv9CEIk1vT4dJVKEZhuEGaXeVHqZ7OEIs8FQjEEsq9eSvp9zppq6HO5jiO8
SsP/FVAOeSdgU4xzTywMzvjvy2wt4IU1gv3iLTkNuQnZkfQkTdwNgJ9N29o25lGR
h5F3EXhkNbWWunN93pzYp6R1DC6UqopaaeSJaFayM3cRSYiVnGHaHX+t7voHDOQy
pUSMiC2iDx2uu2s+8h01QBz9URTqWkial6AEFr0t45N3RxlMZIUhWtR5cT0Rs7XR
bhsk97oOFgiWSC+svFyoeokTiT62fJmtK89BA7L6VP/TzYHETBcdyybz4s4z5Zg8
0IMANO3kT+ECkd++Kbky28MYBYyhbuK66baG/f4NQPN1HJgb38QlE2uqkpAsU4hI
kUJ0bDWNGoPr2kwWCq85LMzNTyWJqR0PCdIS2TivcyEZsYzU9PL584MlfyeLC5KX
uwPuWAMvpQXWzSVNa7QRnfl7YA/nr1GhgpJ0cjRUhrbPTzxZhG6GJa6w2VDMD6YA
Uc1eHgvPSbhFCVXxQ2uu1B/dHwB0B8qT7hqij5c41ayLRAqcvhuweQFtBunQA27u
5U5iQhIFcBqpnI2Dq2d6na0fiJp8wgHxZZqi6pmB/kfVXuzN8RCy28tASUOBfEuJ
/HER731hKWcKkeUl1XjNAtxwTkykQm2w8thoCZgQPe5jLUO4cQAfG2tTXMPqhvMX
RcfKsMlUft5u66ZBVR0Rpvwi0WxQjZP0NcXYsntZ6I8qqRLXKntBb6E/tKWZoR7S
WPIFBUVNlb1Kf8/lyqFaT2zYsM0dH9Tfa8mJ6JcApNh0CpGPiI1csPOjPQYa/dn/
Um/CCtutjS/tViaEOGB6mvRKtcs5MViCZFyXLSbBuPBCQfFYPMGISEWysrSggID4
T1IGH4veOsw5gSiNajMjBpYJuUsi7YWwNxGNEV+ZpzFzLkQta3hHi/JnaIRJHM9s
UEG7IexTCFrEQ0O9YL32F2azjL2KRzbNNaOu6ztwO38UDRHUCxI/1Tzgq04o+Hxl
lXgClBj/z11bsKdLPVNFCz4r0luacTslzOBuLWYqhoD4RNyr0JeaTyBCyYAaqbx6
yOaLcKTjhnusQOMdDe2qJSHON3SNR5hegX0oFUVGu1Uz2nMr3uZgnmo/2vR/LkNt
HmGniisbOZadBTSSVVE1KWwpD9NXwQEYSQNA4iCsOEwtYYxEVz1gMH3EFFiKVzWd
lZKDEoqzBcfI4gJIEkWnk5GklK4YP2w9kRcS4xdb1h4ZrDXZu2i+KQQjeR1BNAne
uJfUW7wIcYZuhjSdgmjO3dRaE9r/EhT+1NTxXZSHRfL5KRVQDvbs7VUCTeRacmMY
VXZhRf3h9cVqmgu9/yDgHIhlGYomB4LBlLmixHpA1ZMORMO+VIxdl0b2nrESa12X
RTmznkZXI9QITPPrffoUjuPQclvIUk4/cjoOkpLU+zucis8Lbbtdduno7f+yD26a
lDBDhIFcEHFGeei/BzpALCsSJHV7kHYkIL4asob8zyM5UDiGFMOZ3Ie1EE1i+I3M
md9jR9uqqAWq6dcxN50+GT9+Mb7Vn09+XYFbmVCc2VNv5RGSNBMd+SJ6mUJqcfLv
VVYhPOzzvW7rCJ2xvtIfbiLwygkiTeXmFlp0see/vagJLeWeKRGrEr3zAZdJIz6u
rg30dRWD9N3dylakImyYnGlqj0kSAYL4EVIhLSzz8qPLWiIv8l75eqBmpHDI/R/6
2QOFPg1FBmqP5sfozAtDh0m0jjVX92TS6AO8ao601zR4aLI+zlU0eFXpMcoxGx8K
ckGAXx5pHYzsLT0vOUwfL0RLUZdO6uedsICg7RyT/Vvi6Fzx5CpKN3k3LXYDjmwW
/2p5c0PPMgiL6jwI1E/zB4FCjiGVUY/wtgUshYLHSUiQtFqDN3SB8O6Y0BXKHyAh
DvMaTycQGnWNb18tYjysQgEExK8OEGJwZ96P+svn3hpquDWEsmBWfJII4x8brWG9
KjbGHsHdqeekOjE/XP9SqfgBgQkRSH3ogTdkrPOgCsKFEjJmIKUmU4g3FIaBB2Ac
XPnTL/Z7pEGSoiPjMAIb1Pi4W7VX1wQ9Y6WNfqUAXJJE/FPLd8C0/Xn5/QIbhUGB
fyMjrqNBCbnUCIbZkC6VQ3e3tUr4CY7un2rpmY/lx0NsQhxOfvSnFipXu0tuhSxc
CzD5+Pxm6e1ZRiH9ZiejE7aJQnt3Y4qnhHEHEVLAHqBecZ2PqBGWR+GGuYBCeCGL
AfVGLh52DUsFWG5dcvUwmTOZXsrjZ+tjvXi9h4bV08MTgT1Wh1p1UGk+CBTg/HZj
dsQ6IAt+4MDvIo/L7gkqhdr9nFUCXvoUOOY1rvAIFUiW7Y5cTa544noO19qUNwXY
CXzD7201KBwBjUoyOD99tiCXNPtmOBmJvf0zKXKtex6ekUimTRhLhTsGOus9HnSJ
5PaQZyjDhOxs7ZzcYgT14s2NdbXVQSQa9vuXP1O67Kfp7Bc52jmUEtTpiX53BPHD
te/1Nx/eogASbOL8NbVoHlrGp4KofbvdNbQIhWWufYtUR12QLzLALLVKI2MIumId
CwklDCLFFJvNqNDNhMIwCOjrnrutxisL0LLsGKAVj+CQwg8cGpMpn1FJz+alhBOn
hJFuDbNDtmRUMCJqBO/2IZl6WtbwlX/cV/j0tpCPXBaxKD+ozuXPNfilpWf/bFt5
HdxxojYa17OfoyuFO95irygrU4+87hlsAOL+em9fTymE02i+q+92BYuDdmY7XnOu
HfHl1SHkcx+1on8cfa8VuoqCaity7QV2+cOR7l9rqPch8HgYrW/1LT6Cb4LM+l+q
MNVfXFnSDkSfuS85EZfZa7IzQYTEDc2GslJMIiU4XvGcbFTVLHFD1DLN5ZP47NC7
tnCD7S0f1CFNuJsq7+2KgbmjeuLO5wf+vpXO/NYxxCV5hSHO7GZQYCsC0hSOrlE+
cvq82zNZQ4ywiQ385z9M60kv8ejZUezItxRJNZHho8BYfS2uNeLaLHwrr12xxXO3
pwGDhDuSTiDgPBdREKhtAXUVzQyl2w1NpzQ5RnBV1Je6eTPJKcQiGm9StwqNntFo
HFdZ0UtUDvIQ+cIIEUltFGoGLsDrMDJ/VEulbz4pB2e1V/8s3XgwcvPZoY4lQHyX
tcWAtuZv0kxRrUtvOFXZ4ovLYRx5DPE+Ng0bBeXt4cCLnA0yK89fQvTby98cnHQd
CjvCRNpl6M+hWvzWo7d4SydSRLvsmJx+ShOIWvLYzo0WOyy3BZ0z35uZu0bt308c
I3lU0hdNBHBSFJ3r+LyDYUbXIQhBVnY9S9aAuVC0gYIulBrL6G5cB6BNISVdHfWB
jpdIf+fVV5N/MydF/Ou5X3RH/xuxa/W35H5Gdn5F/eyChKU0x1FDnmrm8Z+i7Hk4
umZyVQOoy+dQ9FhZRguoy2bR0l6ANbJG2HTCdiLGNco4War1fW6hoJtdU7lYuVi/
JzN65f9ijm7aaorVeIuIVhF/90teObI+0UfHkZhy/lw2fpXcfO8QoRdvfyybIOxS
iACEbPfhvoqv1ZJ3jyL1iIfv5nbqGnufGnJfdzPCGzKHSJN9QHLTHhjP98GgTIdu
4oHcMdiCo/YsXfdkgAXa+mYm0l+a7uM3wqpxs7YtI3pGIWXSBIM9CWdDhJy9PKON
yHEqOArkv7m6OpN4yvaQDNoant8exZ/Dpb4tZCpZU9tbSQDtRYghNzS3ha8CfUpB
8HsDp8gPDf3DvBMhXnL8tcbAn4SwSK6M4t9mTsZY9DVmCkdLqhB7UtgPzn+wnCez
EXg9OFsbLwRX/TbmvPIDJTFypOhMK4YctDm/0TZOG8XMVSO1E1sa56K7kI15TZmm
Veu9bT0iXEmSZhTjCqBqum/5kqF/BFpsLZXUnM3XquzhguSTrnJDC/C1iFdlPBqA
ZITIhka25SKC13OG2rwKxRZ2q9yT6DnSQ4zHSYYyEdYFc9rvcFAn+rMbS9e+bCV9
irY5qlC9z68vh+93mw5J3sXeqZ63PgnI2fFrkpJ0Ync6QHvPwXiCmavBFJEB+j0G
4zGYHKWilKBtKcXjRz9HSIjkhB4pIBqAlmQTKXrY9Vk707iJnNiDTZz6FU3iYAQ6
exK6Vk7lOVa8wLtC74hfWTqsabH4fP72rrmhrBA0o7MZgCJ7Y+IIw+R22HOEBitz
ftqv6RFbqZqMnxmpyU77u1a/si6A7F0O1/yzGLw8pYRB0xOXuI8tzCSCnzhWDHRs
ZR6xWNGbAHKTqJQqBfIwlO1Vlv6RG3tBkcdBAeF3jeD95kuii2qUL/OH+ty9AafQ
H89lj69Zgn8wYJejuVn/820qfOovaXjo2nvx6OX0stXSqJekAeWnmHXx2QdvABSH
XHVC4g4urqlD0FG01hwqvPhSe8KF2x/4pf/dBbcAvg6bL+aKNzalHhnCdsww+ftN
VWfPM97cI7fcniz47tsmGdSuAxDyGSjyJFVegUfbPSf9wYbd4kV/8+Xs8kgy7NOA
400xf4N29FHRfYgbhH1XbaWg57fNHbwC90TOwT9aC9Y5D2rJ6dpge8RqczSQmkGV
mF7DAeAZn9GnuaEFv/UGcYJRpwIX2z3/E3OOWs1O8yxEuG4Hp+qLDjNLAnQSIDHP
mbYneiTSfg6U94YPsyRwYI5o48RX+c810SVqBBrGnlmsnpqDnLGmhdAoEOpM2sEF
+DnANMFkrtOIKlTF6KG9pKr9DWSKopdDGlWvktHComso/YiXHR3BT4lif+DXnNY3
DTNr7kCcGrMwYUvayLk9ME/Hae6QBzCqegi7nV26yEOXPriClVBDMaUbntIb3lWV
dQ4d00XrnS3NMN/UY19+vJ+1NMtmtclPW4kSR8J2TDJTwBqb0xmp4XuxSblGa/LN
a3Voj43VrinHI7uxcbEIMXLvLxq6Ifsp/4XodrxuSRRwGf+HlyerK2/vwvWOgtzQ
aPjvSN2N0OEui9kofKxRBVyjWOvmQVkgJ18ZHKvcM9866oDJbFD2x0oi/NBdzdNh
KMWU6LzpevQTd6whbmqQWS0vK9qUWo9WoP/zPJqW61tHiCCkOEA6D+4ZJXinn9jN
oXKRwOTCp7wIF0Jn2Fm05riI2KCUWfJW0p7uKmZBypQVu8GMrsOBQh1KlhnG9hJw
qhf01/HwPP963VbX9fBhrdL2E1tV+IJh2FqnfNHLdeCEgSqPVrrBupDHfR9R8fnN
V4EuPCvhY9fywVB+C3pnZCwJOHCmq8grrPyLJryRcbaqbdzYdakrXhPCXrYskpJl
cuCZJcu/eCTtiGmJbqpG8aA5gaT0fCWBdYuJnELLUWpXoERF3NbIDiZmAmz0bd8e
ITyEbaIdMYrMqTFmiUhCln4kjnCiDNIzUQDDyhPXBsYpMj2eXs5yvJJi0l+VNlX8
EMQpduxeC8d963eUKJJ4mxB6lcvmdSUQ8+fIYFi77lDi3bi2pz+VhomIRixPWeIm
SKe3jhNdvuV1Bs0uonuSQGC/73UwkOOu03WhXZranzAyYnoW6TKMOU3EGusdip4H
o5Ol2y2YBDHRTm6rRPi5fN4JC+hsHZlvOFR22JPvHyQ6K6Y9TdS28kON8RY7YqhY
qxG8Kpkgk6jxmTKCTZkzZeztkeOS78SL1UfYZzBA01J861HXpye8svPvVwX7unV2
ouj/GqY6weoRaxCASte3SDLn2Cm0UV4jWzpSQNa+ZTCpyQJkKzeYFvhhTm9iaQ1G
u7MdbSSBjLt9K/icnkRKBWX9lDGaipDxpILbRDlwPVi4HTAnspp1Bad6RPng3DhY
qHbP4u2WJM4vVExrWZtt1AkAiUk9nHwarcMKYjam40vlbJp7EzB6OhuRgQ1dn50E
COztFPjb30tdzb8HyAFjBHkg8v0NXlaiwpqjdMN67kOJs2CdA8BrJ5babPKsZ5OY
7VnGlimnvdlVM9qag0IkabTQBD8p5VoURMkHXNLc8fPkMBbPpvi6sdBs/IJG2xME
aQHdmaImYGESD7Z1LtsxLDbTHSNtfxyffrrI6HhOUHdcUGBuWtepeDq53imaNcHk
cxTM5lvgzAi6ZfxdCRjrO4Eiyg9g9o6sbA9Ij3sLGUZWSoXnC/9QIe8lKOjJVjaI
Vl2d8mUFXMiBslnwNBB4FkDQMXxDME6BW13BV3vFo3UrxO7GLKcTY5ipPC98SLQZ
lB8s8XlIShuEqat3TjJVBEsEcCkydyEqep4+fV9/NqK2sf/sIBbQTKgJU5pi56eg
IMmIjPXCHQ9syVzj5Ps6wCAbNqEMBpj/nKmweHV/RjHFYnFX9aqbA6OihrfbFoSE
G/1k68HeJMlucYzxanuv+qs1PVQjVItLsPD0vS6empBqegDA2C0n7iPxEtmHXgPF
SJVqvVXbUdvqDPU91QgXIEDARjjyewAjg7o0UnSBSj39WPuMoCxO6PWiVzTzQYyK
y35ZHlp5KrTk0ngtqGVxCDd+i8xDDJUPgqxj9dXy4sXNcJ+qe3rnDBC1JzeJNoyd
buifNGf5iUK3hXxZY23AW/O3vsu9SuHcZ6u84ur3Od1ihabMhPDi6y5TaHC9cwrQ
HYHDKzh2RD48juB0JGmuP+Ff0ZgsVQ2BAhy7ThODh5gGl93wTMS9AAD9vU0t7Cca
KTnPXRGHu+HkAwIjcTM36y1bO5EbKt64X528IeuNQdC1+aXJ9+HmwQ2PvCgxsj5d
OwwwFoY7GDPYMdmBobScw54zFD5QzISQpHCJbl5UyBTWzhdI/ONLqa79xYodVC54
zu3qAsBsD5XvYl1E5TrQJgwdSgDNwx3hh5gE5c1OWA+K5nyNbqjX1uT7zjeVRI1s
C71tXQygejAVkQcTYPUv9LzGR8WOSBHTe/HUzI2qYbpObuRdiQiWeJ4uAP1NLwFp
IfWQAEiTmmVD3maGgtYL9bKaYEGprwkzT4A2RDtNCCMjfWE9y3EeMx+N4gagZ8QC
AueWOOCPe11MVd2FMssUqsVEWjm0SOX9nxFlonU7GIrInf8LsSSun9StVsCWYXBx
NiFZX8797xeBr42nG6m+KOLTx06AfQ7oDijTMmrAuVu/Gf81oNTuxIXdtsLsWy2V
U1YxZGfDilR5RF577YKkp9s0bNrZcqerFf8t+qSFEEWIvO9NYQc/7pAa1noe5zdh
GPXje6tloR71wjKQL3w+VIXzF+bUUdW2rEnbts6QNjtb4xxYlkxpQRBEnyK/7niF
QMXtqqmuVFWpvAKiB5fWKZDtZF+OmfJCWEoH6Ij2BMYo6ak4R9X0f78phY1P/6pq
p70d8GZsDtJ5x4nVsw7e4E3Cnc6r0QRW+4K+eYWCSN0KO2RbOFZyPo0fxmaL66y4
1POjzaQvN7luG8qeJncKE0aD2r6dGx4f7m/KAad+a+2+heulv40y3D8j0sVYElO+
zOTUJVrdkrbEcd2Ff2BIKu82+ZmliBYBD8a4ZimgTwd33YQpdqfusNIFFRwb5oIs
Soxkys/4TUiBk0DOrJLEKP14V4TQJF6PRyWfaWfqMq2Lmw2G5P2C5Z7+yqjubcp3
qFoyZdRnvFIouEcxIBLMJq0gTzzwquKTkTbr9zr/mDkzrPa1QRX1gb4kgnOnp5bR
UeVShT57AeHY6b1l/ue9pEdXfYsAdqA4iCSDo5Mb0Ebj+Ia43zH+BBqKIco3/U0x
Ds5THbLIbPLuhM2HhnN7BlbAar7/k3VnzeousOjXFlTTnKyqgco2Zrc2G3xIAWXU
JGOpgtUVYgQ0j59fGrTXbh2en+qBQpCY3tH6ADGZKt7TZm0u3ST0nxhHS3U/emuI
yzoYm1z/aTniGVXiiW166EWwdqy00NOUHMf08RtleTJ2iEmn4QGMyVB9Y8sVpyj/
qE2EPWVhF7DujSZwSfwt/swmEj8anadpWCAvdMsqlRMSgEjAc7UpfRTBJuq2xa7g
J8u3GGUys3GwzOrEL/tbiT3Ri23/pbDXn4bdZHwWvuX5dzaAXAse24FpheJEflFd
/wRLaSTaFcMHUE1m0QK9fSqnI8XO42DLomYSNMX/kiQwT0nozntEKqsCi0oifNjm
7RLyAZGzOKEjj/00i6An4WRvNXIE25s2JXfKSj0O9fPvy4NbyGuFrgDNKx84NMf2
ov1q67tFSs6Gkl4Ysn90rcXXSu0rJZEP7sPDI2HwZH4nCaXKfg7rBLv00mkvHDJe
qN1qW3ApBc0bgIjmyevxq+Z/5uXmIUTe/BsnEYKZfkx8wD38oZFeMp/zYjWO0JU1
tWD2UqcBPh3VFmo56ljvEmRHxeM/4DfEWY3JPi5tXsJG0FUumAkeIsudPLyOZ5tb
FIys5kfWmy3Q5hWXuz7yys2iNW429WCFbVfceJ92p1tjMM3FO5Vv1I8gEvULXgRX
0qJG3LV5IIE4UyEvsZ7MMJLFtsFg6xoS0iSt4vjPMnYmf9zQwTlaBOVxao3Ql3iO
+rCr7qVUlzB8g7LKNN9E2SC9ydRmj2VNMzCehLQoyFyTOmUO6Hv6HvG2c5eqjOXT
WhHBx1tYb1KKY+9/96vf9fGx5HoPdxwI3t5KORBmULEIRxkMONgXu5mO2nfqVVfB
ejcATtq6GQ9MVqvC0UxOjsLhNt99WBgd8zaZDM75Igo51mX6z+PNdmGbLGe8CfUx
TOV8oKfA71wNREZU5c2bLq0AgtRTcdl9pwlTjqQQKNT/5pSfhJNQwBZo2NUsTRgN
sAjL873Kb9sN16RKmuksQSbBUJs+q9kovJsWnRLBpkiGbT6evYJ6KU2GdOzxliNE
xW+dx9zBirzEG7gBkvOy5M2VFAhIVsz1Gyr4FcHCC3fXqLslHQDqkGEclcMwZsAc
afGiyZXFPb0zEPhmewOj9HhLeZZRNPBMyZxlkZd+U94fx7dlpk1JvUbAAyyeMreK
PzTdKz00JJppPFLy9t6RvnwaMU60Hr+nfINO4TxyJZKajBZLgyJqHq3GWB2M2O7D
XRJ3FPYlEMmjTZmalx2qOILVbMq8dUmxirIEvG7hiHoAZeOAh2wvBvRDoUK8B/SA
L07dz3F9SOrPIr8xCU+BphDADQ60/r3MICf9VB0jSICAGbhCcdwDe4aSuPfiKao0
7l43tUwvUPDtAKyYZB6eQFUFMsMiKmLg1u4k6Srm+wWJZy2GWYTvRw4Xn3nz1fMh
z6VZ1w++wWul1gIJQSCA0dHija4tnBtQeXx/hjEV0tMqN+xQXW4RBg84b/q5h75e
JYJpn60jm0mN1CfJOQe6FneOzKnZ5C3NuT8DgLT+aa0BOLAru/8I3iIGfFOIipUT
yTy8gTBN1jvw+yWx7SoRr6JW6Wyk7PrbYjCNp7KikMRb6rVRBnBw8pwsXREromQV
6V5nmx/KOmGuc83vlzrHg87NMTnFOqGDRY0H7WANi05erlCGUlxV6EGAGi16Jvs0
gRlmuTXzo9Rn2FNeDORlTsEJxZjQb3TMCDmFV4efN5skFEs0V/odLUc++GwNzrno
wM8r+hziGqJ45yNRM8GElY7A7DfQMI5LYIvQ1aUw3lUbJLPfHx7qnUPI+Ynu6XI8
RqUinhKT4N3irLq1SZ+YkjbTGoXpzCd3SRCejAP0MqQ6HNM66SDxdWNA/JQxR6Ff
iSpGYJFT2en7iBhLPapDYpXxnPSsmMUmfT5IpkNPY8pCLtzL8qLp/OZpsMop/XvT
wgm9/sWpZghAlhnUyVx6QEvj7Sl51Mb3xLaqpTSKR6R4RsIzBO28XQrSgo0EKG1U
wRwgWfti5uWwf4PGe42nqZu+DyihvwTJlqQsvRKo+V/eVE/IFLqB9Le11gFWxh+B
8Nm1iGm2hdMRHtORWqU+jDE/7UjHCEXD6SEqvTuQO/MuDw7UHCFSpWBgCyWZCSh3
OZFHTrpvLuuIGwpavAiWHBWuwfQi3t7rbA7XMzqBpmRJmKxz4V2cxVpLkAofPi7F
7UCka03f25/B6rog2c72yLIBz7WZV+RWCcj3ehvNB4LwUxpoMIP+wConA9PkeE+r
VNjPWnnY1TYDge9s0aiwrmeTS8nUWprQFoRTHR8yXbyI+CuLqRlMm5PhxlO+GjxC
S0d+n6kxo3gvidbvQUIC95v8IeC0YRYC1cRJ7prbxkFPuWh8pM0NyUmLRhc3SHQP
4BE0L/QGzh+dvwoB6xGzS+eW2vKuSS8+TbpdysoAfeO+AG4pQq3kQieTl7YhfrRH
GrafWPdnM4cmE++SksR7ozKVdCXYFTX/j0Et7Ju8lLxKldFjgOZ4hZCT8zbIWMSQ
1eLyv9VEBIMO4kMD3gpyVEbEQHPY0hrH+FsunfNTvlFUH11EQ3T4k284RKN2a7bR
41h9gK3nwaavxX6cGNitSkTA2LDEeRjR6K5QiitEmUHb93l3OSLPTo4sX1CH546h
BvWUoyiiqoyVVwmRELgbCxs9rtV2wz/CaFgE1m3lyivMHZG33bNZcibgYGHyUSvc
35hO9Wczetbp9O/2JOpGv8dDH2T/o5yByzZcf/Rh2I7iDoXawyIzZPIdIQb2nebw
WhaeqBsE0lyU3D3ZCLqNNoTogT9fjOgrJKRL4aaoi3FdO0o4AsPMrrd/9emPVn3c
oJV4P9td+jEA6X1PGfr5od/be9/9KndL1PHvtVlyy0dl8Ka97wNqgFQORWLIhgC+
k3L5xSUsKD1tAx9OHUtshdUMW8bu4lBhQB7RfewgJvz8Fjpc0Ch9wsKdIqYBeRCf
RAbJ9psCN5FCVlOzYVLrjzkA7LIcbgsO3iKc5SOfNUdqoaJ1JZfUZfQGk+Eivebw
ufLGgSP7IYOS40fz902S9TqL+p2HYnfrmbwxwStyYb2JAGK/QuX76bEaX8/V9uLn
vMNJ3G9kaFN1vyhH6/bcvjtYilDV9f9VLVp5o64Rw94cNuKRTHcoJKzMsp8AT3hd
nueeaFJ5f3JzURLa8dkoh9u4qosT6OsFSTOseEzTYuBin1Iy/HKVbHsEQOkOUphN
M0YnbVvLxqFzYcnSQimQskFSe4Uv3Xs2tIEsXN5/DEnY8iv+piTYP0aszXvCtEeB
wyzg9HUV4Q9/4EFY375OuYNrMJQB6mi0LuPYixiutOXgPwqBzQGDHfIIWKSSeahW
dti6KpQBWtpd5f/hXBHXKZqDhMQjUygwZvyrSkAGJj0N6KJUx0n5ynxDHpL0OnPs
ecWQE7EPHdpMIVuf+AhXEE/+w9arF/7hkMuEY9/fLARTsJRENlKau2I97tRPUKI7
ubytMoTC+gIanqxw2UmpEunY0JPLvpQY7aiLO83yk4plm3tnQ43swhJh8lSz9iJW
PnKhcO3mMGH50lQkgMvpwmFNNw9y9bMAuwxXvRKVkES7uWADwldVN9jNn9xxxK3B
QjX0/m6fhANlTZmXGgGBV72jMLv5EST2B8WtFPxFPUjZlaXQOdiUn5Fw6gmutPgu
FJZyhnl5F+GAB2TsrzET5h76YVZzBgshy3rtMyuMI34to7Hbgvy1CoqOEdndj11X
ZAvXHJmiLOyhWEbFj2cW2Z8azTpQ7UEYOEH41pnzgw0SOyt02D1RLB3BLZt5HO88
xYqgqqtnO3LgFObybMLBmeepV3RSy+baFRa5FbU/A8qsb2eVW7oDhBfpWI10r0lN
Yygiv9Q3ZIM6YWBjPCbpoL/OUA9HFyIZ8A5WjFdHB1pqeKKIqsJVGRjt1Iq/8eUr
uh2rvcgbvW393Ikj4BcB3ow1MPUnSu/ERROknzFbaUykKlWCKNSDG0+B1fu2BEcr
GNOCsZX4LFwbBCargpV7wIMg+w7K3ruO/YcVgS9ne/RBPg+F86p2yTUGUlcmEOnj
8WMLxo3pvyMk8DlqqOP218xAYwUrxSkyEGTgQEeuYhjPKL6qz6go3CUsFvVSJlO/
Akg+BKVxrOxkA+20R9fykW1H76dQWwLhEGLFSMTOaKmAa16lEwoG5075ZuvF+chO
a1jfpYK96fzhzIydZ41LVeATSNUMX/8+Tp/kA/UItiRYh/NVV4v+TmiKGrwe0LT7
W6x3LdFHuVFzhWghx+POWrGkBw2rkXK81JbP5cP+8NMtmLu/ZEeQDrEQbQiRtH76
6ME+5bfLLn6JOhbC/sDY/A4Zo/S37fRHC+RJk7O2ckfS058dY23oEU/whBM1MrSm
oCzVCc0lrJMZqtHJwGtcVgcqyF3aXYYMh+qjHP41uihYTwr+mAHXP1HJEOtvXmoF
RDxpSGAgWhtLIsACQSmINqcOBdT/VBNdWbvkylFo0WfexWb8vWx/Gk+/PAP7vg8R
XqPFyVqfZ6k0d8daGVNmvrxRGFhZye+2xt43pOke++nHtiAvhwAs5FCLrVdLaFV8
KToIttobnLMTOkvXlCAKZoNUFeIL8keXwtk8ZibNyDO3n4i9lfj+HN4WqtPgkDE6
248hBvhONqWCY+31K0AzzEBR31nMZ/+wZxdwsuexKc4AyEO20jmHef+qiFLbL7Bd
23nd8bxGyazW9iLvlAKzmn36f5GIWxhMXtlJG63x7+Cg8szcK0S38PJ9A1++tnj8
+TyZwLg7/8Lb0kSUHzVNLcQGf24gsJ1C6HaMbCsM3Jsj1xyfbQ2RSRTTTLlGQDXJ
KXFWY7A3oPGrbjtEXVfrREP/p7QSp2jdhkmXuXlS0NtBfR9D9yRSiE0ZFjqxAlRb
MIXrj+FBOCcz3CLlvKCpklriMhA5ER1zVmpnIuW8gQcfoTklVdVoctMpjhZAL6lU
WO2ZBhm7WTaN8zg46AgcritHpzOgqzpIvbRJadaYks7OEM40OhI+O7AQHPxeVrTW
zB22bGJHFzJDDLqg8o5D+jmQOx2hbiq9mM9u+ZDY6EAN/KHceQIaePb4Si3wSqGo
JCvWWo4Pc+tlG0IlIe6n0RrUEld/54emO7yvXFZR3KwEZ56UFLpMi6z6Xd16TYq+
dLctptq51G6C/d6ZMC3YJLOU44QKAn8cNTNKMtlmVRM0jQ3TstKGtIu5QNHjj0Ic
IilqrlLGQ3tpND9vtwaYwxJLwW5m2FrQ8EIel6X1buE6QpxMegdJnm68oAnwL3QO
wSVIlsBhWFIQ2u0ff/FI1kmmnKKr+CeRArHNymtqq29cgZhhrYrz+2I/3n2mSdVX
jf2KA0U1/RDiwq9dawQlAo1yKZwxUJGKJOnmgZGoKsQgKeQ4pz5Qi1zGACe9eaV1
1xuwgb/SJ7GEzcpevQoO1DNchxDW4QgJIbRpfer/3cwC/4Mbz5UOspHDn4+tmmK/
+hkeBvjFdYg6iX8/GYNdp+EY5dYRw8ypDurnwpcBNkPZWzlH8mOisErZzAJ/PL90
2WJKVLV/CaY3dlK75aJALgObX7AE/+OTtwxwNTSDxIKt5AU5r150xx64ilDzgSFg
/2KB7MYTAMKfLwbao8omTf9Fc56YVnxN9Nw/iS82JMNUstMA9AsnGh7B5c4obMRN
i6lQ+zeA/zvnZwJgjmPkzaimoGSQs7u/GQTPnVeo92jjsZkQZ2Fa9m4VF2vjy2Vs
E0NjP//rJaYvtBQnmsPpU3cQ2p9tHEmSMwDws14/CsQ0M3CW5Q42AhvmhudV6cEo
JskUhZgf36OaCjOfXrWFD2BqIu//D/2RkZPFTKbfUhlWWKHzyANDBsofkV2giInS
1ZL5sLaMRl+PPDj2EI1taxoJ/+fS7pxhKYRnXAXesSF7Yz6+Uq/Mz8Wp3Xjx8n6T
4zutAHzD68amDIbk/z6gXBgw5HVC31DDkSFO+gPq0xlZRiPeKxRaqxboOIyh/PX1
MgenAEzvHXJlWMd78lnTE7r+P27aRczqa+9A9Xzm6zL3rCN7DTmLtRaocw2gru4F
GSzMJf7NPZRoqsto87Tc5BHVACzUiHFEkJO9CdpMBl9FbIzzOdx+dq75XiIzkjyg
ZXL3f1YCwhAs11A9nLFA41nYQt4/8mVgZ1wpg5+o6jmw/jyLBxj1zImAW/Ylk9zZ
MxwQqiuUirhrk+n5w8j6ZdRbJguE44x7kkWh+1nx8OKNwkuMC+fDgeKDSYC1eIj+
Ufe1KpH8WkP2IUCx1IXzdxEnsjTa3N4/tccvXB5TPe4nyzHy0GBQ0N9LANReaQNE
tFiExi7bBlCRuH8mvOYKf2KyGiABZN2m/5QhXU1t2IjN7ilRQdBnNTi4MZBr4Jhe
4fvrk2uJoX6ghwDeMifBJPYaKTYFO9B4VuJSZwHeR0CjHsmenESv70F4i9M/oGpF
perOeNOpBj4NjnihaZNAUszJ5QhCeKd9dY2m/iNBdqi48dZcqWhfuUm7rU9zfFWc
rrFIH/GM2jpDWg8iVnVYHC3/qOID1Zqevk7XKARIMjCp0w2+jITIpXmZk44qAdMj
GYh6mrIIq3tnXL96sAWriYpa2BQEGPjneFxvYi4A7EwtMix6XxaMpA/w5ySl3dDx
lkTDNMaq6v7GN5YiVeTiWWnUYnQoeYqMCVrtw/g6t4Vy7KMmduyLVkqX4xJ79AUy
9lo26SHXUCyme1Kj8otM0dH6MsuJqjmY/ZohGkzwIdPV6gXaF+j+VecXiSIwXn6y
oHbtP0E+HKZgJOb1H5u0zlEWjbB14RMUh+Kvr3RYG8r7Y1vJlAM+lNBqNKfZ7YLD
WI9WXkxZQoXqS5xOxcUxc9Bog6A3GpkrB5XJ1tWL4v8/jQg0wbXiSynGiHQWLR+j
cuseuVgkbsUD8fHRNmcp4MnvYp9iQ5mF5PIczseAm3wns2tWGfsDONwdEYUvlh2b
XmaYBK6+KS8SYtz7BDJTRHT4Ffyy2ChNd9s0pnaA54dODIakvy0xOTc6T3rVf5hf
7pSXM6YNNISApWiPEld9QWxTdKHdqkwrkXrDGm4zBp8Xlz4d2ByoOWpyr09+QsCu
gIAaxvcMBL0oxvZyIgZ7gAZwhzDiqETcXVw2+pns2B+izMOt7TmfggRrUWqvmirX
0swRYU0+X1ggIyWJ5B8JSNXY9lefe58nJrPqjvNjoQbs7sFV8gT6stjXL7MFM57v
O2UpKPlYHVzJ9rBT6UsyJMd/dS/ybfliu/BjISmePFJtCnr5EvlhN/v/EXY2Toq2
bdzf5EBXO1OCfgbqEMAv0xakkwMXkFRWgUjuGwIxVupcY21r8yW5sxCuu+D8aCVu
gzRKr/rvUhEntzwtFIfO8AMeNeBuLV46Vd/+WL61tXHh14HV9ult0GpkW8M5qUwb
oMN216s+IovPeb84tjbH6F0xIAhw0TiODNyuTgvpwG+ZnoOBPf/SSRDa/4wA7FS4
70M/9PZi6I62xei1a8Ktws/Tozr3q8NcMAG+ma7CZnec74MNBThK22yWKrLwH/9c
Us6TBnDqu3YdVOM0hh3zsb46F30mUO1RDO/+4xG7ESjI4jFiOQlByjWksAW/aAvy
QbMOg+PKYNRubQYvHQvqQvsSpwF82EZQ8XuhLu5XIFedELvK6pAAvS2EHahlsxR9
/VvQwa/T/+7mb782oZYQuErrfpqlbHU0lQxOJTHr6PaRVbnRDhaGKown8OwcQ8Xc
FO5Nk2GcA0i9fsJY3955c35AtAFRWLuYouUlqsC69BzupCSrQNMhNIuMG/GFHQo4
HGYiAqs7It2dgcSdRivVE8Uoas58bVE+IDtd8eEsiMJD9gUXJaexPycQS3HMdRBf
vXxerCFDfLtcbrlDFcGTuy9ohfKHj/1XceCJrwlYh/fhLeQmZQqFLof8y1H9cIgq
9cESB8pSJGmE2vbz2gTd5orOwi4gF8cA7zAF0uKLwxY+wTV/ZestygwIqWUvDm5Y
N9FLUy9S7JH7WzPqHvPyS9rVYImmCHROyAD7dBa/Zmou6SiIfP7ELLNJr7ANHZsI
4bHAYoffxxbwM1YHREDKo8vuoHPMSLn2H/CTzEFk0CQXrnpzhwEfRF/w/B+J+x0x
2QF/uQKZkGmJI+ETbW2X6205AqdHbVu8gndcCcafATyHBuC+IHHJ0bPR66PfCYHG
7Ig9MXS3qjq+aLF13YlH6c8pbix+rwXbROPPo/+xtafDTl+4PM+JrDbdjRMRPZ8w
dH91sECQNonbjchhx8r2tInSwFvPyHsu+LPhjsjFmqBeO7quVXvZAoScp7mCYGwn
kOyoRd15FFpXFuD7vAm9PfLEpyzOIEqJ0UnjeyiUY9Fs3uE4iX9okac/uvgI7B2o
nuvjnmcYsd2Aa7AAjwaILAF2BrBrHltcP1a+uaAxxZmJPCw8h+9FvGf8ouy5zxzM
nb4pJsCmIbDiz2FVOrwfptBf6WKFGCSK3qyPDFnuXkGGfl5NxrytiITmQIGqIpv0
A8Lvfc3Ee9FOkvISQZXAMV0VAb4SZ4aTZfFDPLYjZBinaWmKPchWe1f08bWra12L
bZ1ggKgO4Wptqwea6uw6g9hTFO+Nn+/Pfx2tJXojhfIW07rzBl1XAOK1B3p1d8qW
sFi2LhOI1e43I1xryiVqvHZP1p1hgPDOrEKqWrX9IDyNC+q1n90Sprs9vKffC98V
IDzeJecSO6LFhp384CRZFhqVJ9Bd0pLiIm8oWvv5mZhWTaipVLTLkiW1wVN5Yqo/
FaPfCY60iBq/cjqcTDvvBPNsqiVH9t9nKvnd4wh8beYzQ3QKAeZgnf93bTZPJPnd
pbSvmDjVHpK736RfH9SCL6IrQixg5z5Zzw9KQW6g0R7t06F/1cFBi7gOIK2n5P9/
f0v+4AGjegcf+pxGKvIs74U1qBrfVnwITd3jRbyuXqnAd+VWA3sdn8eAxlICa+0g
a2p5B2I2M96fnVwWyWYIop5V1Q9kQ2xNSvzkuXjE8kMGtycAvz0EkP6Lv8RaGtHt
+Q/G6rHlX+4HXAiN12LdQWqhxI1FWgvyR3QldDkkXZWDOgAy32biIGtF1ZzS9Jmr
MRNDADjrSUd1A6v1nMay1Ddu2YWA3vXJ9kZ6kRrm+U2KAcflaGQgkKXECUDDRT3L
m61wS87YqPOZ5G81tCD+Gow0LBwdaIWNBPp1vTcXVgtl3sDd3WT1dk1Z6x5ZyKYO
bYXj0jOSASV4cO5eOcUCM7q/RKYqHVDDw6RrGFKyMfvv0fO+nCkl5AlVdOGsnVS1
Bj5geIhdW+RsspgSmjAWjo8vK9BNObsRjBPxzJqJqTdzfAfyAMCtjo+PzCgY5c7y
JSp60I60RNrEFgMWvjrfhrjdJ9M9Ae1g6f8AOes5sVA2YFsCKRlodmW+ANVb8dHB
+REr4/Id9okxZI23ITHrpfGdfJXXUZTVzRg3DUDx5eSGdQPQD2QMrDrZOKkS1HUC
Ru1r9qLeHCEqkETWNGm+4q4eqC5dvYwo69tIsggEBW2NFSZBjNi0qAyZREWfcpqj
sHdwedy3fOsMQ65bWO8n4brZ+IewqI3U5cZ0811AiBpZ8x+iaFo2FIUvvsL2ZfAO
NU3wfQK8tdiDuCDrcrt+bq7MZ9oeVuP+YOfTZ4lUqLHMMn5WeNe9/Rn6O9JbMEvE
z6H1YfKqad9Sa9FqtXl7xv6VdOYXxAT2Vr3iaZYrVGKk4xHo+b8pZP3I0mkc4HUx
6S9IYtU0RSCOKmVqP7kimh87nvvtVxtzZc8ozC3qy1s2/w+07CR86c/njzS9U6rY
9CYrcV6JJioHCLQDokuvaV3JVtPgpQzy9sEsTzcbdN0FNNpPZzQZrNQyLeddFyVg
SRsgameqmwLXXqqRfBz7Cx6SB+teUI8HbuvlPKNVyfCdpvXU2k/6uBj3Mcd6EJnc
QNp6kBvMXWpZPBm7fb4Bbmai2w1IXeQgxen2RTN95UDjV6zflY529Z0cqt48bmrF
DG3aNa9KKOYAhuDHmC3Z8/AcwGKWj5sQhSJ/wQWHxan48l6UxYHdWzioiSXlOwwe
luJqVDjIlJ/p4wHEphV9kZjqi1EjHS5ATQatAS7NYEE/+JIR4+e1PtjuHsVMIVk3
kOE/shXwGlyoDuDICPGnqvt3zR4rXWh00gmB4SZItZC0axdXAv1PP1j/edpJJYCk
v+zREsZsE6HDAvYLm/JIKMSV2JgDkT6ulVL39oB34rzDROZHG5YXkey9QKt1zmzu
8CQKQcPy2GLuvksqou3xqHTB45dAO+sTHnrgwsjrRlEGkDLvv+tVjjVAba0P4ilH
iViqHwUbBMlZFUN3r9IqssUUx2oaHwIuHtLznQu//vXl9e41rMAHPOwN0p/X2mj1
TIynAtW1cnf6Z4+utEJtxOWghS9TAgJ93Dkx1o+hHRSKTkyJCYV+8nwjJg7icrud
c1w/24GpL3FXBIms502WIPhypl+o0AmzEqvVzDB2yP42HXYi5/9ffAqZbBQCE0Gr
ZjYrJ8Is0v0ZHcyr+9NcrK/vzTsocT3p4qYLd7kWfBgnJooNpkiAsY5Q0B6SQ/ER
grDK3lr7bCYdLQ+YwldPhjxRgTRHcZIx/0ZIezmkk2NkiG0dNfeYqrqXrKwmZy7c
mZcVjqwint+gLIGab2oqKLM/dfVcp+8fPQSD1qUCEchU5E3cgCDZ9cRG1zheKF5N
uRTgC/q8kF0UxUXCICSWjk5Ax9Q7eMWtkCBCs/t7RipCwdqlN41bJXDVl3C+tpaw
6yeGFchD2ORA+lvieJTMtGmZAiv0NDlnyAmiire9EebQpbkDKlc2dGgXTTWX1yJk
DWQInIQ/c3rSn390w6btJEpUhSLAX1Wm6C1hcj15vcwsCwAkeskaFrChYppeZ42c
MSOJipjyTvNBd7pH+gx7xX15wj+h3XgcUHuPhkwMp37uM0ftGpfn0D4HtdstVNY9
z11NNVwgJWIaRLJ9EuY9okKY4kGYrE4KtHr/7+Nu3+xQ6be4SA1yxq+xDNYJS9/t
LCwnXJ2fobcY0GOXlD2up5h9gCNNRfu9IgNDcleKh9vTj3qDXVi4uVFaIRhHmtwP
sX7co6fKx27xtqLFhImKncoBwdS+1bwSuQsD0VceWnXpxZOOB+etaSwi5UJYXinW
eS+2zH7gU/r7V48NYbaSLNloLMVwBQTZCIosIEY12Eh7/oqeZLixjvxHE1LZkBXX
yESPbHWR8xoClKq8Wra67ZWi2lFYZK2Xy30wXjydAHIz1v3o5lO3kJbUpp+GBjTb
tS5dDyDExUQ96xb5nCfCPJMMwjDURFzBgRd0uLdHsFR25DDdtvZZ3pPwvWVcOtBE
dEsfm7jW3T9kOf6dQ0XixAF2MB/2waYCcnUjDZwhdQxhnue6CjjT9Idi8dliyWjF
xxhE5iq+hyi7Mj7IUvB9HVg1Pmb9krKPG6/xfa1XNsdheF5vRKvnRXYRd4Lmnyms
HNsW7YkbHaNryqlsCvbKCVUquKkUrYGA5uv9S87h2XYE45G2z6Rm56soqGYwgZ1Y
yg53vyoKKQKp5ttrxwtdTLB1PE5mx0X3tJXbDD713eefPe24K2SvJqRLHogn68XC
jspOlqy7P9Tt1Gk2WasQ+azB7RPd/2CWpkU2teFqMaKmY0vmaB83VaIh9GAu+W+U
LUVzqx779Pjn6G35JkzscIW3SV/p99Gt1VuI4F4QrekFOq+On/e8GLoXigqFULvn
oSg9baRpzTQ8A9qjpPCrDjzdqDOVxCkv310Rv4e07rlWmuOhFqFhqqUZADXizic3
MZbnDoaMlmOzyHaOTt8TAjfQahNFeeAHUt6iJiSIOhez8z68Flo5eKrwRLTecAP3
eD1YD+dpEmtqg8dVQnO4dZiyd5CeFpGbPfhuOuIXTU5fK5JBwi/ehdRFHBFIPXfs
pc+WogspIxL3XDkkHXG9qjBrVs9zEooquV6joQMhRZVA9KY630QcbsZ3zhkG6SYR
n6TMghrm+5wviWZnMUJ/xz/4xJkcyS3xyRXJM0SzMug46tea2WE8rTlpKyWioOHq
aPVQVysfcjUqj5v+u13LHwvdd7IXTkaEjMXz2HUgX4AaeOsI6E3A9rHf/hyvlZJQ
a9TW5/WkJ1LPtgmjM/kw/8pqWKX4V/Ch+l1+ka4Cm+eYtdnQkZJbaNXY0jAi4VMM
m5CJD5bpw5FmEpPryyjcR7lLLOVzFFe2ILaBCyl1M0lGI3bjGYKSvfSXhjgo6mIk
oiTmT8GnUgfnk8BEHAQm9vM0w4jDHk+OBXZYGDP9BuJHwFu327F1Urn1uGN6TRh5
Z099lvviaQCI5BEJChXoaCstiF5BLlZSKBY5hPcGDztu3i0iPTySjBIx9vMwUYIR
0WL+DwXYpOx+4RW0jra5hMPFqfo1+DxaG3RlONp2h4LEgWqUDMc4qH6JwBAS3Wh7
dLmFmO2UomHqWkENyLp3pB+KbesG7gs+IVvGPcPa10X/Ve3dKbpDNEvneAm0NTqg
jN58tOby9vIap+uZlg/YIzZaJnRh0zllFQa0B57gNI5yqKnvKMRrn/cUFhFsOg6E
cikaIo/sheWilfF5VsK7uZZquFaDoNSYrV0wN47Z06c4sog0xIXsp51F7WnItZvi
yZWVddIAHMOwdvotsH1umIBR87hSqUjIkVMdZ8NKSdt0xe+i7uS2FETZ1tP8NRsw
bt9N/O8WW/yPs5vTwHETv5dOANm6bpyMVvUS/paw2b1A7ieOsHltUbiTgwY/hawF
CceN5g6CUlvD+y6FB/pBjBEmfTpXWu6wBfSPyj6OL0DYsPdnQhTdlxfcE5B4bVPF
OeXyVaBK3gePUCarjOyvTWK7AvcQBVToTfKGybWV/QhJQydybaVqcl7IO2vWHJ3o
O0jCmDc4kkcnSMXJcWbCrnwg36+ocnTG/28txQ/AFRt9lzyUbottdE9wlIiquIhC
257rpHurw4cSREZKoyVsIOWpyv55pG+pHhYkv4PFiX60G4UaAPZoAvCFAT3QkPHB
3t1sDoelb4unSdH9etGQBTWjjdpT+icKUdoHgUkDVTHiCZMhFxQQIB+wHgQ53A7z
q2yF6Vc6czA/jWxnxOAw2UmXpe/8/GMzmHHNZtBXN8C8itKrVhtfc6we7oUdW5lu
mwqn/kjN9fCFQFLDhWesaYQZIAtE9NexZgnStP49NAKI7bxxyk+ZfwJXddHlPDJ6
zOwxP+/9RKSJ8CbNc0dbLVulvbiy+J1UB2Qq6no28e96+RkcRXoqDye8ss79jANd
WdnaiNFljnPz2gfawA+YD6to3zuSCaz9ZbK3A89OYoayqTkrBZEzjE9QEOA+/UiA
O5fLlKLyq3QiCUI/+NFzfIG1y4op37Br6JMrl/7++VE7RTmR3bTfRRdOLBkc2DTV
JjzFf307NzdFCh9BCIWoYEa0QL8pdxdwNVlYgEZrdP+Ko24B8cbvlCn1hAouGRSX
f6kaW7NOUKna7WNK+e5x4HdMckSKh2ezx8kMEjyktiRbHtMBuMlSgXHXoAw0Unsg
24AqQgpu2y57M2ZhrBLXKg4THbk8Z37vueDmRnFv/+vuQsDjQ2nZDHw83fFVh8fW
L19uwdV3z6kitJAo9dYl6gTSRiOVsddC7G3rNkvkf7Ss84L50NEPQJ8VcqVcGZs5
p3ba4lwPzLejCfGYlht6/XpL7b1MwgYxweKsGgIhLJ/CD3PnqlrEQ1slaxVvOKJJ
Xlw+gqBmUFwkXoAC6yN55P2Kr/DaNoNIOxDwhhX7S9GK8+f6H3Z/yALLbgiYHYvx
qrwqZybcNfWKQvmHtqEUkErh4TmHNE8mi4/rF2aEOjkOXdC31TsqfG3aACxIBNoE
sAkQhk3vHNgktMVR0slFEYNdQ+Y6wn7OQ0eX9+6ty2E+flEDUEQgarHLYb1jI+dd
VTbp5yIouP3dYo7tf28oTlOSaTJJWdw/B7GORZivg0zDLMOag8xtPMIopZuKlhdk
QGLrRtCftHcW1ICA1ZjcO+ISOkfAAQnWXFR/prgwzLtPrOK+txQsWcyUHprx4Tcj
TY0FqGvE4XZKdF6YC16sybhZwUzSE9FFzPtsQwnO+nMXBmZAOft4k+I/x8TlKeCq
98vAKA8SOpRAy8YTXgK9HJWxWzIR2knBaYsqA/9x1yG/8VeYLGN9KXpLolxWpO7v
MpPXz86BYtXwbYvFyG/EbosrilOK/vLEWX/gPSH/8RVX9+P/ZW12daeeAAdEARF6
a/qjANbCR2bO07ttDbz+GHWU8QHGNY928VDwdmjkCDL8VDLF6sGo4NsX7g6xcwit
qBcH38+kFVOpsMC6msjdCqEXR6Dzq62y85NoSeon1OrFxZKStT8+JVvYk4TVLTMo
Y+JNcpkY89ErfOB8vN3NSXO1mFY1u2Yy9S2WBrH8d1j8W5A8HxQYD8+ztEKSzfKw
gaB5z9vx4u6YD4EXXED8fBAng9ArEuNxf0NDmPZlKd7X7QqzrCpSIY/e3Gecml1K
55Zxl2OJQDyAhXwwt7QU2mJGLYLVqhJLSpjRyvNQQrWgH4Bk4QdNC72YP6ZcG7kR
oQhytgW+fgqo1f6bbqDQhJuniTqJJsjrEyzdTsTYPnsgJs7ySlsl04IoFlFVM72P
e1lUW5xBRfm+ndd4DztMP5CQOooBWjjKTm/9Qxrog0u8necQQsKcIpW0asriWe9g
PsUo5a0EKTTo3i2+x3+UPdOVwB3vnIWR8y1VgNAEYvOIWihwpqeTuIj85DmWbwGu
RKFQ7SXpEQviL+/sDyqQRxOVsKixMcp3DNWX4mbYgHkpebOTzh5XvyALZhth2yhA
WPTKGWF5ZAT7qMomO/jYRUqJBWRq0YCF8E5AGmdhvKNTKjWvEZah1benBJ0pChzV
VjDDJOf1YvJ67GjBusWolCe6roBKCUE4b+drJ/MMnqKmoA/kxcmx3WFzHJh1Kt4C
csQUTQP9YVYJRs3GDwImQ0wUBQJChRMi3zdfVmtHA1Rp4vDqmdge7ITFnlu6n+iQ
HLY6GeIWUnFHphcLUUwAprHjLlAfwoROqMBx8GQMTzR1VgHWPelK6gJ4RCCTtARF
Zd3rtD/KPtsGeVhDtrxXBZwP2acRaOdxLK+gKKpLw8LvSc8UQxs3VA+XHjS0TjU+
cHKw4bzxqzLqyF/SaqkkiW+KxyaX+/8Rms0rYrCurkYJQgw0Oxc15PHIgXQcVEeZ
dmv/4URTuaUJllFqfBbEkYA7T36DgDCc/ELzFvq8smHlDayLeYyJ6hwFJZoe+xef
OtotQnaQFB9VSuODXpe9e/NZ/V0ikh9Yx95ZLQFikbURtUih27CgFiMGgT6hbezc
AJUyXIDr9S/Wxr5MKsVV8gqD4PIgoV/GBy1oSSr6sAwI0AHtprJaU+bdGYKJDUPA
He2yWb610CnVeTN26RrY5edwGAldJ12fqJW9BRD4Yd2LvCHagCzuvIcr44CUWDh1
NxeijEoCgQmScKqADz2txReCF1Nq4LWUBLlYr4EXi3hPy8lYz1mAr0wzIIW0yjPt
t3XUlJPFoNP9YttiwXqGr/BSZ4ERkGJAKcR3QRCVnHkYeXLK18Es6BBGLcWLCyKJ
/AlYRml8lIQI9yrNsTk7fOuwoARPuRK7Oz6oX/v0sNAxU9ylnNOy7/RJ852Ip6zS
TDBHDvL2yFMRvHpVo3i2hANvq3mn3QRc5bZhY035a3VBAc5PIgyfjTBp4JYl1MRB
ynywSmIqm49BPYaSLoNAKg5uPx6hDqtSX7qJ2G9XqanMtG6VlNTdZUiBoedKZbzS
peVykN4lo9H9ZnP2KRpD8bb+LBjLx8VL42j7zvvJelKSCy0tV2r7SQfM6zDeRkS8
HroHBoR9t6mrGR/8pNk0xJ0MP5IT8SVQ7z/LlnRt65TsVEmf2SKFRyo1V/It5pFH
OgRZkYA6eggqiHP5BidNnOay+SxIDiggkqLyioVI4+ZjugdX588tKkGMRxoS1mcG
9eb4HyDvD6extHCVr0LtkSLsy/hY8fGOWNGj+ZUG47T6CH4YYU0TRg8ykcIYydkA
2y+RuMP4KFbxJq4eKm3pIM+t92wh4OM10Yk1zlt+xRKs0T7vuJFNbnFqtIpcwRW2
FEhjJV4YBsUwx8wDmcOGQwR7pYsfN6YH1vU4uvgdosLL7wh26HDJZNR4maR9jkEN
SqXbRIzHmPed80O+LuDCK8IgBDPhM/XgF5KVIXXOX6ED/SRQoeRtXAjaKcfw1ylo
o4QfKo/sNS2gmDMRSCh7OATj16qGDHKvuyeoEp7UCfVs5dJuHovMRGjUO+MPwDNL
HlBXehUgBS5+GF6dG2tC+NDVqNqSeOWq+PEv40EelrX0YGfkIZ6eadJFbMG1AQli
IiOklB41bmt/7/w5H3b68JaPcMhk26T14mdWU+yH8AxOtUV6+MU7NEZpBzyvHpiS
2qV65rRVA0Tx9ZmGnF4JVxqV5rUei1DCZiqnsMT7cCcAYZoui4Ysd3oo9MxJ4L0h
eag22bm7DHidOS0WNt6eHu757omYxNfpJGzKVv15ru+gm5IGM/KHXVspnu21HkLM
yh18uq56oBFiDv6h5o2e5MzXMTgy9D63RRcR32tseS7TbQcpYN9t5xP5mSwe9DlE
GPikziYpE8NE0EFlX4J+DCjMzigcV4WkMZ3b2XXQnOaJMbFHG/fl91mIcpabnDo2
yg7fI5tVHQP+h9mKGtelN13lgzlIi5eAkCkIUwGY8lWheFD3Le226KG4DZkH1rmx
BDJS+DiD5MdWu1l9Ng5Totqw15D3P1T503oLiJ3j9e5W+Yf91U+iuu7YPKAXAcmy
UJLYmN+HB0I2DPhj3dc4cr2fhd10A2dmJdmggZqHTQK4wH41tuApcbwHRWEjoi4y
1bYwDbPhYEIxsmorWZQt9Snohg0/WsqssTsH3uomWIEKNsaPJe8vG3SLRPOfWf9h
nxobTKqRaXl0wMFTJnASVTsoCssBmVoQiAtX+ShC6vMg6t0wVSVqaivGg5+nGOuy
qkoEN22wMGt5nhIoo3TiJ38lygxhO2fSmyClebrFIEDMWpSIp/HAnf3kxuEXHeiT
kGA5fsi2rs6OH74Ufqw3rYJdouCPsNh4gFp9pTc71qmA+AY8kAzCRB5RvOVhebj5
4kWxWksYz6rmvIFBlzcOPR+3ZnSCrwQHqBOjdSI3WevM8Z4wpwUqMPG+6lzMgZDC
ydjJG2r9W11aG6n+vYi0llwRioLLhkgONtdTPPyeqDIAzMf7a5emd4jAeayGZBqU
YK6wimw/rmvxWb8Lg87eYufGIiDG5OUIgevPeMp1cxb1K6Ez5ieSAMkAYln9v0P6
5zlgajhxi3v+SY18KH3/mj8vb0heG85lhLrkjX61vDMc2nJNcHymYV49ImVxfK6C
U2glquSdPxspBrIcnGq151TnNRhv/vdHHwqEfU1+gxbqnUCunaCNXeejm32owEBq
IXT3TUnh2OxRjSZNDw/PCCSJrsl4MzDe5CDJ3dGNBuo/zTXKtBQEJFgy0gUTvT0/
Uje/Ti4XfiM0yjZIoBBJoevoUi+yZ9W5SiY14h2J8wenuf1IJN9RRp6wLjgmYnUB
oYo97b9H/jgLIvUXGho+sZACL6cOsxyxgmI4nfGx/r+NbCWNO9iUv/0G3FoHtOAD
w+UenRjeW42hW3V7w0u8DNXOVGtXp7K0vsJYfT3l88rH/rhDBd5O5NF0j9GDJSd2
/ruZI8I4sLnywBb17giPEOVUIYuYiNFoIw1HegUsqayXsW8x4ZCYQdLJTPAtCZqw
4IC1Ms8GI4pjZJU6Xo96GQcsl0XSGqkftTFwcgHkM6muYO4l9WNLy47Z2lxNgiPO
HJT5BE0ec/4Ow12TC0UIQi7lX3+Qw6RK8fwawzUdK4DTui/dHofvnq6bjEBVUObn
M5P0ISlERzeCLvOBkhPYV7oZSeRdW/eRXQ90TXRN3LL3ZNHbe2V44TAo2cXPepYn
+JJLWEo1PC4zLa8ffCyWeUlIB6wzoHw94AjnBF3wNOepKIcIzQjNiHMRcRlHkWaD
/q/07HEzYO0HeBD6n+sKk+5QqJOO9ZwCswDUg28daPkf2bu7ZLHqLN3a8Ewa36tW
8dFB1DugY7N0I17U9kAaM3zwu2K3F/REMielyO8qsMi/+6NZoOYKb96nDX+cNcpR
wYIsICklYV4hrLEgGQisJNsr+uyphSyiYhIbzSrk9xU1BX+xigwkuF5qknZ1KZdB
ualT1CnBUYCAntaTPLF+P3XpjB6lpog4ODXzE9wXUvQ1o1o5bqkdYzX92XVM9zzp
poDDjbYJGeXiq5CjbYyaSBTDHiWJ51SUgEcOquIztNP4B2bPQzuduDwyBsdLuxV/
c3Wcj1SgGcYhGyaSbvTiiOTkrBAXzVfenKTbPaA8VyFLfSL2kU1m0DZEwi+fi3YB
I8hIQxankTtRYgnyXUVRTDEDrpB8HgM308veYnf0DSM7mXisV+Y+m96LvaD+V7AE
9t7LF3I4ebzGb7O90lUJGZHO6zicVcBsNFYZ761coyJqB0ke9NfvSsGUD011g7AU
pSXkZnLX3hEsLmB4Om9o3TkAjlJzkw3vwJboIPqOur3Fgum6GVpUE5VdOfLXkdWt
8Z3X/+7e5qbSAGNv2diITmpcfrM6s5bJ1eWx16JX/2zFJcfAKgI3hy2z59D7FTUT
hNhhCSube+qYQOV4Xh318xF3QvOM0xGYKV5KMLq/4PQmmtYsoZXkvG3t+vdbnRt1
+86pgWrzW4mn6H4CmbMNzkufoAgNkxWspIumpj/qMaQJZ+G4fUtmp1ZJmaITOLxv
yL+uFhDGsQcSKETuAZxaC1laoNGXKpiRSpttEDSAKyHbaLabXXix5DCdxOrVExBS
6cHnB7jM7erTFsiVNN3XxAC/iwA24xrM96w83xNmOxBq+Rn7j6HHX3qXNW6gez/J
qs23tcbJ4nfTtTp1V8gvvisQZQ7F7BjrTk4yZ07P+EAY+u6yL2At/KOvEbLi4Obt
M4FzgDO7UBI9QF2SfYeMuOJtbEQ93xqr4ufSshrPIiKIcSujBz8sPK9P1ZEQn7bR
6VnFtpVWhQfrdXg2T2vOAMcRgbEuKdicUkL+WZydq87s08slnu421mxAE0xuVu+l
ahHjhsw3IkYaYTRUkvOhiQgbQT/gBv43lMLv0iA9OOjvq6yjy26c1UYEJYg99lab
BUtTsj6dthBNy7o+K/AmrWPXE1gWZg0MigJjPQl5ytIkwGKWjaSMArlxUyOC1dve
GGVcCFi0da4MSd2mO4mkzewg44qzy4m7h16kmJhBJCCBamGjAXW5qfL+lWuG41bE
QjoHfhZ+MUyvjTlgVGuJI41L86Ng5cLDhhyB+yed/twpJ3sZCGXImBFVSxmCAzXq
sbcicziRC9CKLVLRzSh6JbxmG0UokRQ8JqRqfgvUut61v1QVsgVkvWnaOnWqUImq
c5JFL3XTsjG3AVrGDurByAvk9uOyw2xXfChSSSMNNie3LSyboOTD6U3NltQi7nU/
l6rHcK/PHV3MbKVUak+qIi83I1zkDdR335vKcv2Fe4qTQuprqDT+8yGkfBkKy5Qk
iOLM9DeC2/NXzEyCGPrjEG7w6dGD1fOQT2yyYk5Iu4AMuWPxLrC5TGdM+2gFtGQR
M1yqTMUuERqx8k8wlG+BNo/YInu2BiBmeaCkj+XLUT1OridFA0MjVHDmTUku9ioM
tJrSl7hfVnMQnwxXKTpmIjmPeI4UvRngnF1CAThU0X+IocUXJO86GYXUV8QgqbLs
GlbGRVxxv1XD933wnLQbGi/gS/onZJxw/FZIMZ+zqAIaOgu+Pv86ttWG/kpcEonM
EBInvk5ldOCVv054cRgo9p535H8rAoYgnPYCGxlvLtxtbryIj5/mddgFbCkubwS7
PZPAEjsFRqfvcTfCj1NOSRI9u6Our/3Iq/PXT4pAqOCkaQdO3a/0DsWy2g7Ppge4
eCTZtuhVpJ70cBJLlW0UPF96LUPqOL/EOucMzjibdlJf6UzrDSriQKbbwqFuGVUA
PX9XSLyvIVK/46D3aWp9G/7RtKEo6kvTefTby81Ni48tZc4qgEGdlaKY7NYEEDdq
tJuZSo3DRY6pXsL3GFNDhDH/Mek0DOhv79Khp8z6VMjrbZ1cRpX0jVm0BWZEX1nz
zMVe0O5q+PkpUwCd7YFJAPxrkNiEA2mU+btvvFHLlO/fCk4OAOMMoOlXBBRlONje
o3/MemHEsfSkD+ItdcMNrhX0UpF4b09OolunMFKtNVQv+8ZwdKY2Gx80Yh5r3hfL
KKyRd4m3caG/mzfAeW9IwYTGVFs0dajFv8NxbvA0g+xHKJb1uc46oB4J7wSp6EUL
aTiLMk1865GpW9KrFBoWGbEeTjOB5WnC7UcGeiF3hIw7rZBMmN8EA8JgPBsn0YGW
476JW9c75f/ED1pAlSwID+6soMVOD2tuaU6nQ/mdGyOE79+ctncbXOu9//iX7toY
OPd1nUiNttlUgR5ClKnqiU1/vZJ/rxMvq88Yyh+3G8PKsR+I1hjvDdjOw2aCCfM9
miBJRg1GwYUsSa9Fx6bNPM2SYVS/3Lh8LwdnoP2mLhOnd1SGTcohnWPDT4CDeGjq
RPUzt8ostp2/BIPx5D0aZxLbKhhWD8C5Uz4cOzJ8oCEZsIkU6AC7nJGZHuZt7aQ5
pP70fdaUNIWxX6LigQOfQsuhJoMyH7EN/KElj8cQ7TXA2CSpwdKTzZGY8F59d/li
19LvzYksnpCNbVzeixywiGaFpjWebRxWJWKAsjPTRprDXek9oLHr5t1XUG1X4SF6
FFalL+c736uNWzmPTxetxPxI5QOCbYQWkR7Qbq5M00j5FQ9GD6PcYV4CNtf6/eN3
uIfP4+Ak9+RNiYz2+bwbzPesC0VPItQxU0nMCr18+hZXkHX2GnxJhL3ExU7BEufA
wDp6eVyYtPEyk2mww4WLDwOhrixATLHZDkhb1JohuI/Yv/kPw6uTbvGGMSBakQmQ
L9yPqIme73qEOFSdTQipGKtP4mBqKO9c4AMt7FLJa9PJmX85AvbWRSJgbcmnatlo
Kw6/TdojwuUkopC9fjzl7lmw+BCN2yackdLwxuKuJm7N56lGyR5oe/Yqm/xMqNJT
72VXybdURK4k6V45W0fXckh/qeCZwrKpZlWdrWDiPjxyYeh8fVnC+vPuX3xpkKsI
zfk/X08HLoWuK7s/oM+W9RBdxSed2KIhVL5fLkj4FotNdMxvtGZdChv77I6r83XF
wydN1I0jYAmlT6m5eIVDlfBjxXJx6Qu+YxNFkwMF3MYiFmmQohiSrnTfHFumS7Wk
MnubvmeOGPmYQBqRHfsgRnip2pW/2EB/6WNLgs/0/DnjHA8JvnM20Wc7jp5U9nF5
5FcULPWtVpJiJUFa98XTAWtqkKoO2e370UHusFTU7YQMv92+YmpFreYXkuSBtlFK
i3LdAiCNX7xiBK63SnEFA14Amw1jyBiuOGy4fHeYqhbBZNJdV58e8n35sFiatOU6
yQwIGmHz5chCwJYvkZFqPSHA/a5VcK/IqlOwiid4Ro7/qBriYAv74ti64e3oalPn
vblFFXE9+VmJTQN0u+9HQiRMGirDhey5i8u/EWdZdlD95F5laTkGz9dVb9tlWLFb
ZImzM1wTUKrcJSMUVSlBRgPKzFCKDLoUG8NEsZN8lTvqXF73kQpdIepau8CSsGJg
e1AvQ0oTVsjwrjXPQ0ckeDz/hMRHPyl4hvurvuKDHQjnpPDuYMi3DGwTZThVta8/
esTIeP5OHwDozUnW67uJOoCJrOmWoDCEBxhTEyr6HMfJWtNjGgYJ7sJAHRWepkpF
soR3DMRZcGWF+7HN3eaFc6MdqRmbbTm88FCndVIdeJDtTdmlKDgoPKhf4TZKWhZb
DOHCQbtzA41LJd4WdlQ+Hkt2P9JhA08Pi2a3TPOYHqDO7UdNBuROoTdR2Y1G//op
RNJ+soY8U98K73VLFEWgbbn3YEFufiUqcAFurf+wVL8FMsp93c9Q03gKkf81GvO2
9dez7LxUzjnZ7yUcDGn8MCQUyYZTsdUnNTDdc+rp6Nt3UInom+Zw3Uip3N9FO0Xn
hdZ6C+ACYpUnAeMn2oi/w0dTaJx2JbZXe731mSs2Z/9Z8IRaLTITcdij2Q1+MlkQ
ci0jkoo417jGZu24VRAgpqt7wR1i55C9Tkhh8glMuaZ+KPENxt7HQFWU/VpItMVV
eMsjzaOY4C2eWBN2N5oHpSctx7JMgUK/0qPUnn5XgghkuiIyX2K7XB+lu0irSSMA
eRpiRSymkmvAoz0dHpaY0Tia5diYy1TPXtrm+yG5pfRiJKfKKaDlQc4s4xlpnx8q
L3jER35+8RErNG7y6D1fdue9U09FzXyfH9KPAJkqJPQHVkbUWAjQChiRHiGCI5iu
vMDS4+slTmSimjEaRy5xeInIHbqUxWjmplUUSzxTpEwpNYjb5+FRT9Dj6NLXOab4
Eut627csSv5ogboL+MX8DxPdCghgRierlQtvxi8ErURJIRg3unAqetnj2cvzHCWt
LL7gNjA5rqI/Me6dSRTuyLcNSaKRvxElmpJviBH0VECIn66/V/cK66uJJU0smGSb
l7SijJKz+MHM+UQZmugoizZo+6S82dPXC5veNsnkjCUUyHvPjUM25TuLfovvodS9
mOcUzXW6BE+ZQmtUUaT9fJmuxoMLWbwKjqm9sp9gkJL67TFrpIgq8fqsDCp7ufq/
0BG1r/GPA357UXv5btu1pU2sIhi08rozJ+romZvJZy3RVG9v6pDkza761hyocfAm
AsZQ0ceDAAHIVU9qbcc0wA/KAWQ7IszIfoDmpxhbteiOxML40H7rVnCdH4nLOAPs
/2GGdHDgJ7YIDMX8pxPtq3yjvLPYHRWFQERNAWsoUk6pe7CxK8cy/6C/eiLVhbK7
dxBfI03IZzGJeVgWgFsXDQwm9YyW9qKans7Ev8Od6iYR8m1Yj8yUcaW1dKhupxtR
++W89P/RE2UfSh0NH/eg1mhvXpCbHR9wPx1uKBTC3JOY4swPUxOtRIhYFylXa/KJ
epTyQpw8FmZ8pln3aImIr6TodCAeYOSVRm4zy1cRznjHRQgCaEIBF2iWvdLK+eHY
pNb9oOV5gYIUCsimNP9zPvzgDmX7y+BGKt0R698g/NGeIcbwhnyKVqD1PoaVZ3tD
tIctflGXZlQx9GRaV7QybDqOYH6HKC0sPipkxcv7xZ0P4nOpqr9e9BdPCdpHNYQZ
o5dL8Xr/nur4uglj4uoli5s6X0k7/hJ2L+m5S3YNgLCOEt31mhTEBt1U0JDm4MgA
CKV6fvFZYH+OEj507WDtfBfjK82vwA3uviic6M8jaCXtI8ZuwwOK57Ijw1Mc8dAn
Kh2sNUu8m3geBxlwyHZPSxrNmUq9mDMOJqTCDlOG83i2nPafXQ7Th8dKTeyLHMzo
5OhB68T3bDZYLnF10H/zBMnLFENCCvb2G0D+AW7TE4bitLg7bhpF62jjxa3ZY+2S
S7ZkZH5voCcLF7Wfm94oWsZS8hnU0y2tkQ6UvXsnhuIe4+r7+rfiZEAjBCm7skUU
YPAZZKipwRQ1qIO56hmLWC1WNMvUsHM828DZ/9QCaRUmVwEIcM9bZZcOikb4dH6Z
SisI1CHZnnxbNTkR+fOMEW85Ej7KMdi063nkMQc3T6hfDgFsX2plo/TiIBRoZOnt
4DU+3VjesJVmjwOm9alvgyO8cg38KkKfrqeOXA1xwWkf6/QnzzCyuSvLTHPsnr3i
HqrXogp5T1X+QtqvNHxYJXck3sD8RESvlFyLXF7PzvpsNGGrUPenXK8IylTqsHbS
VpzXLVpKRNF7H6qc8IOKLO9cDHA9RUYOjZdIBjeyaY8lCEYjx9SsXIc8GK1Yndy0
eZd07FZtmgseC9Jkz8fkT+h7j8r/S1gD3QEWuXorvpyJjeYMIzwPXnw+X66qvkG/
q17Ar3k2xWJq7bXg7N2YM4t3oLeeZZVM0rQAsDKBF1SXzOhtoaIDcm+Y70gVmc9+
Huc2yXtEmIFFFPQI18aNiwYQP7dWyQQLHSa0Rrx1pOAQ5NNsRzvahin6J1rdrd+x
aBOiY6a6HUFAo9rVGQTAAXZ1ROv0GTD9QoiYAy8kis+OZ4im4ZynPpq1nF0YYdEy
Mc2fw/m4vnY8D34BvMGa245U7Cb9PU1wsjt9dCv4JprnhZqSqEus8F5cKEGPnRKU
xYh9VPBggASMPMN6Tiefe+q2pkDKklvUqUyLniFe2zIEAZnW+Raj4jzBS01p0IeQ
y4/hzc3MKmrXVTNgKvoPS1KDrV9X1e8GbPpl7VXQ/TB3zZJc5gY59kD2vPEmXvd0
U+wRq4d/PpxVSwoMTng9FgKXgE6F+Mxe5r3MLI9LbqjZd8jDNdCS5KOEVRgZ8fpG
Pt+XPRr6PynBObjMcSNCWnWXwo01Y27Y0jFNW6yY3r+SY4ozyCffau1t1vkcfjxE
C0tNaNXMZdt+ArXgKHoqAs/hrDICKDKMY3OJRqfD6lE5PfqsYrle5bIz+AfRCI9k
Slni3nULXvtfpHr9SM8TjIfJQ4fBFtOmb9Qm737mSkLSfKS7qg8wEAYDv8iixHnp
veRN6HX2zmpVR3yxLqzAaV2mysT8K7uDCEmuosseqiWMAsSfYYYa683xjI5uwae9
x0kMMuxhmNUKTWtyVEyiXp8AeRKL0Z2kMOrZhnJth2QvFjc0ZYNnOg61Uao6mg0k
U3Mn0MswVoTxU2KlPrZV3Ws4JVWUBbCiSxlZlrIC2TZ0UXhP9YG73UKveBL1pG1D
sBfVm0bYynpTHsrgHrLtLphTRSvHMs5vBJBooumShsZoiCzrk0ukuHPAnmJVUohV
0o8zUg6X0JzT0XiB0uf9ISAnjWGijhw3kJ0siYx6fXP7P19xJPGGToPrWCrSDxvp
9IwuNmocnnIj2AqxXcFf0/2ri7r0Qu3uQsH3CbSR65y7UVKpy/jUCq1gvws8lBWZ
9xwuHgkf9XIVWDJhQ5DcNo7NIh/wcNSvCjKg7qLCMg2nhr6vr3bUvIdad4TEU5Aw
iMBxj5Gz27Wng2b4Q8daPmowAmYkbig6mJPDJ+dQiQt0SxMf16EofEI9PFlIRqHD
iz/KoN07E8x/ZHdTaLBEPxGUpNLxpE3TPokkc9RmWRwiajMmKsbA6H4P3+Nex5S8
3OXAEeEF9DTq2G7lA3ycd+tCWm3tKIN4d5jKQ5zcefzwE6WKY10ZPDmzW4N6pXRR
DU5eP5aqbuiKyZowpvc4/BUjjsyHl6H7qYmcGFVHA8ai6VCPC9DGA7LP7PrkddpU
/fyBTYg7yNa6JfvQ7zXLwckRmCpUeBXem1+EbM5ZkvHIw4oafF+vqNWGpL6Z9iK5
izcvv7w8PUob5YYzvMHjf3nF1UFvKRrrctL5iuaqU/45qGercAXZ1sxPdYxQFK9W
XiucdfyqLmR3c3NiUfcKRXwM49kcxo/+Q1U3Ftg8mxqszsCOUB6KCLqn2frE4gPx
qRVwy/j2jFQ8aEyX3LVLrPV9sNy1BSpaduviGw7BrHnDvcSZ/BJAIkuoShxSbTuh
QobhDcCDkDAdwE+GuehP6hlgnhhJKQ2SWRfZLOrE/Qu9PZXnijU2S7kNcg5WFYBH
dxa0yL891J3HpOOnUQOXmHN3orynrXel/oaT23GKUI109ZOb+gQ7LhTq3ZtX1WOl
iXw1B39bLm+oszrg7HD3GtkSeoEPEa8ddClOzM4ZORtiPJt4E0Y5ecgWyuKxflQg
PWksspjmHJtA+7xFAQnNOEa1MAG5yR4A2/uC0gkoILUhyJfObYQixkgehOKvdaRD
MhoxHGdtVw+wtq6ZCv4rduxV65HiQSzLmpG4B0SQ2APV5n7eTOym7/AHTwAFRNrh
NOKXhw0fFwH3PuHLnqFVFQHaTwZJ2JZM1PORqY6yVGCfl5SqzsevpPC7ywr1MtkN
QRC9nr0v6EZOEwTAQOJOyrdi3exQjkb5XzQoMp6gJmue2IRqLKENuT4I7l2t8GPQ
29b13rYiggiVkdHvFtAieoYl/f2jFoLgmlU6Krf9YbAYgyZ6RqoNlZDXSXEYa3pO
JDRNuaqbe+EYt8LHWIhrix303KGmuwQ55uPYVvOxwpgDEWuai8QwUMEqRc236XvI
4jlSmPcIcXH37vvXvJt9d8jbcBsPsLiyvHiqCZ6uMffimqT9h5ZmCaqG4hPeycdr
RBp4VyPnABvVP7u3HDlhV2Ff85D1HUMQbnuOJOCedo8FnPNdKtmMmIDLNeTgHoaa
1f0k4Ev0lRu8oLgU4v3/V3ekeSUsNouPG5b5L2Ia9gyde/O8l8xtq3dHjz+2kf8n
2nRVkSa0B4YGpRlpo212lLCWbeLi8hVLCCVHr5bKa+dzoehj6cT4Esr1xr002dCx
WgRzLSN6sgAF+c/q2ezCcJ2YBg00CdG71dfRQMH/G6sjLbnLAym6e5MO4Tljjl6/
KibOIipP2nSkX9tXMSElMBYoFawTTofAKkn/I6402Pa9zrUkmKgXa4I4kzQcAtW5
Gd2407ZwY9V1msMZl9frto64etGtu4pD56rM+aj7vjodNb/ReAHJHT6bf+2KXvxt
hHAtqezIlMjjwTQ+wMr8mxZkXIcHjB0gD2E84m7iG/9vEbn0Q+c6UVDI3p6Wy424
M3+nJmZEDB6j6jD/269PrQG6QWSXRT6LnFRGbeQ1Qtlu3MrhjLfYGKcWpLyGGwL/
lMnegcuBUEULCdqVWathX9rDxmiCrjIsNCOdHleBPSlX7ROeiqDu+6upp4R3lKNu
WIvu/ZIapMv5SKo73TqHD+URPqUZghp4OJUc08Xwbj4gF5tg2cOwIy7sRBXNYSl4
oPaqtvvo/XPfsXOmr6PN8eWH2+T9JC30px1u+rQSOsOYYlu2Rr99hofwme8IvDVM
YRHGaHcJJKeD2hseGIvzsfjN8YDDUnN/A1olh3yE0swM3ETD2UYwShBKPpzrdLjQ
iwh64RJ+OdvvnhOaxYfE3yXFn1VtdDHi0tsm7mYJW64VGo581HkNsfLr8qTxkYgU
tLPYNjqUIW2D/ARFSLl0L1AD7kUPP5DEHKgHbkdTwQi98+JCBt9knpjNVIjoDoKJ
acNaddDU+RMP+YEEKVOXIB9iEYuLNtp5t5b+tuWFGyjcv3yyHKmcalP7kr5GWMrf
O9DJCNz6bmQiaflldB/GWiG/bN2FfThuL+UX6tFNH3B6aIL8HSr5x4xck5W2OU15
8Ch9njgyJIUWIg1wl9K/SS3hRsDXO43MskXKLGHFrGNQWM9LC2Dd1Eq9xaAjKNRD
QLVPmsIZQePhcI8jB5OFAQKUB1RRPJKKzD5hBq+QRwEAyjv3jao6Yv16kVO0Rmz5
l8Sg9iRkBfUZ9MPCx5NkQrwCFwg77ei6JNBJ7dvArE+cTH6NOqTVhewSuuHZEIZF
Sp1o0kAMhs83U//awDozrWicIkAZ44fn9bxtmZjr2gcaVK6rNCYmft9c5PPigQI/
3RtatLh5Ym+2mPXcWXL/shcB5SvYQ+lfv56+ESf5NigH2UBdSIrF/JTK0YQ0KDOw
GRLhZcPyLszQOGfnqLV/sEAdEsRQnb1sh5nxlLuSYNEI4Q13Swbvs6fqveBnaSzW
zLwTQmnRAVKvtxWBE2+0eLNC+TKwoVF8m/F4Kgy1BaXbr/8aVt81ywkDEW+ygGC5
TrPALokGorg2YPIuT8R1NQJ/SX95pofi77d7zSy2H2Q7mj4jGbSfs6y6C48IXnSr
bGz6lcKuuevbtMFsIN89mKjB+PTkEoCILVLyZBiHCDq9WAmX+b5DEmATKFtTT5fz
NwSvUEKw2EkMOUGRkOLfZenSnZV8oyjPv+HR7TgFCJIDxR6dis5oUqgTzlTbO1Dn
64bYchuGBzSQcqfS4Vf7lKrGXZbxqUyXfOevo4B3RW3uLsZ+IGAI5hyhnlM2osZH
P8qcuVS4gtKNZTyGeeiFTOXCTA7TwCu+nNqCtYfdp1tVnmsWUSInWyuieh7fjvP8
iUlkGf6Xf76AlHe/1rwK4O7uXKw0Cl3NNpOTmqWXUKMKuoxxvVOInI16Yk3f21Yt
eSwFcraFpU4L2TurzA/9FtUerwOUyRgqGxuP20VunB34vvuYHSJC4hDk73aW61kf
sci9T58Z55lgdN3sn3/ANxknz+dB20l6Ljh1q9n4Sm47HSBWbBGJ484e3FvV7bOD
6GmkEAMD5usOIsV56e4+VudMaEYjPEuNgZ2PKVK6ExAax0dZfqXN1att72ShkmDe
Q+CPrIgAtfIQCujJrK4V/5VuWnnWPcQyVes+JohjVxJriv6tJ8juCxNE56kRpWHJ
mX91WBtWjMWj/V0CUIGly1fYzpNo2o6k9s2ew+IQGTzt2PutcCSBeNntPniC979t
km12/shhklOBzTjwt6i4Y8a4pNLd9a8OklWVl2AJNd2wJjKU2lhACWh5tWe9QddG
etzGt8au6lErAgW5kf52WDmn9/iGwwvVsef71n3Oji7renX/baYO+3M4S1MosoW9
JPx88ZjqC9eEBDJQn6bVrvJ9/djO5Xl0zLfjYffwnMyLDiyk8/5NYpMSD+Ksfobb
wJer/djvNjDNqUdjsukwOiJP6xR5+1kzIaVVZZUyYiM+lx4aMImoXcRGv0H8TWHy
s0nx/9lGHq0JzwHwZWM96hbHKGMAHfRt5RzfzUYWoNqTYSKa2a4t+Hvp1mqL2d5A
+DzrhRPLHBxIpKnW00cQkEr2sLFPK3pzMRm51t1vyU2if81W21Mjat8z4MrSFOlC
ruQXDmo+sx2UKH44AUS+4ZjdDYpPEWLJWOhBXomSS3Ezx1Rngw3d7LNE6azvx3Ul
du3JwLwtzm9tRPojw1HwskbnxIvKJcoxOh7OjOnn9HuzB/DWgKs1AXEbm9T/Katf
kHQr2X++mmwckTxRssTEYhlJEPl87sJU+Tp47QFElQHKrap9ZZMGKzlmFHlvJbl2
Xf7FrAUrrGy5IdedS2d2k0I0Ioc0Yf6JKQj8DHmJqSDwW7ClieHxAZ1RUrlKoYqV
51jYTUzSVPqA1sEYcfYDtbvqmHgoZ3E27xtCPUzrNH6n4xkyhpPVhRkaEzIEgT4d
9uezz/7xUSSkNoixHqRWBL0ZDtuRU/Tfs1zB0bzoczaPuNzqEJt5GxzlPABtGbSP
gRQ9VtwGlr9JZMNru8Cq4ku4vLtFCR9E6HKVphSljuyEa6YkiIJXtk3PeTwW96H6
63f0MClYShmccO2EX8vhzDxLNxfRK/PbWFc+fGlgknDnYYFceoW5I3rTMzrM3nJ2
qETqewR96Z84fG4yW7fgGe1lndM0/rCTkroKNc4VqD5qu9LA5POczmOZrHbFTyGs
zg05GIZQ/AdmV7J69JqxiObwmD4yFa9DrQ/PuN6fS6I0zzxmfK/M4iFlhdlkyeFB
qcLBRGRUD5YU7Bp9OmHAeSeigfNqqySMQ/WirBRPAAPWMK7v4kxLHqCbfNJIHzrE
0hY76UkmjKWnLipkGJI/QFDoYyPhg4lLOyOX7Qo0mcceubj4N1frPrxiWTzsQLYh
jhQ/e4gj3nqJdbUMWtVQlpHeb8Gsbv3wR2ruPDX/5sX7LciRhnzXwhNAEc3/plTy
wl+hNjQoMdtzbPepGaDELTai63DSkCtMlVz8S2nDcXfptV9K93nIoBRB6O5x9ghq
9lBOI/Y7JKjcU+zODNd2/najJ58hooO62wt1QPfl+bEHW4QsamwzTbPv4cu8rUSj
vJRwUIWxnrTcTsq4QE6PQEq8sA/lTzcuRHWRpWlZ75YQYFWqWf4rCovLi1bk/+MH
eqIw6yc7NuP7Z6EAqPs++lNyHQkifjZQGVaVr5Aj6BqHd6rrCPRZwDWo5zhR58b1
2XCR1XlCGGk+TgrWo+ycnuAI5TZvLG1p0j7z+v/BQlj2+tAaS51exGmudpGrvDdi
QDnSJeFEWYGzZ9Bct7RY5CCu4pby+F3g0lAq2kEBzkXNNc203fFDPTbM/zjwa7V1
KmVAn+fiVwUmifBES07L6+8axFOHtc+PMZDpzWHyu7003E5tZnXTBu1UCFw8UcSe
XVNg2ZZAszB8RHGtKXlc5fIJP4b9HIHV46ys7leOlMGmaseE2volIuJkKiXVk0nE
kgM/5sDFBMaf7k9dMmcmW6hO//Fb93OgHId8JqLPNJ+EzfDQNnQj6wqeMlZCn5QU
SAdmvJF1bw9a2AC+TLjcuV49X9w3peX9ur6PIDva5iOeixV5zHrtIEw+UsZiMtce
w+k7DCSv4sSA8hxP9t0YCVjwvvrl6We2NBQ8gwlq5MVtnvSsXZqUTnezib6BOFlC
Gct0zH4pcwCa35RRiF/U/m94jdHgzheIKsx8bLeLK6m8b/CzD/im8TSiKrQAY5SI
8IrVOj6QSpNftNOJUn5jc0ld6Y22h38KIkX1F2nM0VqFK/v+YdINnJOcDO4xAYDR
naF3tZ1tXoA4BPmbsiknfoPVGySqLdjJ311J85Szd5Cq3pjqqTTE5348XJwR0XaJ
A3D11FjC0vtWMB/whFROudo0hgSToH9MFsS2vFJXCkzZlM3md6pFOfmfZLe83hLQ
pM0l7pj2k7PWSCRGkqlAPeUOMuDNjJIL9oPOEjNWSftJzEskt9xhAfrTmko78WLb
OGL3tyVi4c/lGEGzRTXJzRdlM9zWRkgKGOFLs0ixwWAsxUAkaJSUoVuKA0RNy9n8
BPYTMj/ydsqWH2oj7/k3SWsTj1qvPMKvj/xsEQuQvoss7sZSQaJSKZ3mcoccsz3U
Q0EuFpGC0IQhQxtxGK6jsA3eLIbqgTSNnODOAkrCLX+BareFVR6C64vXnvicX/mo
g1NJAFswGERX3lnTkova/hL1CCL1yoHgUehV6MaNb4nLn6aMeVIWXb4oHEu+h4CS
TMG84S92tJz4usZZeUObq06WBOEfQF93dzjVUUxF3PmYXIwsvs5xI6XMcevktRj3
utU8PBz+nDoshN5Mo2M/pxNfhdFRFQhoQbx2x5F7xlu0WPKGXM6c6EbiLwcDD6wg
dNojiYI1XzDJIwvRfqDP2ev99qb6ghdn9ikgwbNZ0NqFbSw9yJ+B1R9IgPH0udYF
jXvdJTqqfl7s/FvrwCvSg1dvzOguCKWZ6iKFTIdfehs4Mk5yvMuf5YwhFIcEfVqv
oUwSMPyLH57kQaUeNGMGRTUh3vTJbvC0NKIneQwkUre1SQ8gRQeAwoU9vZjTHzda
0oTea8jOcPiVV3cXt9RvBDEdHTX+7weIHAnyzQkOe5cZ3wwSl9eOfUNJC+vQ0wMQ
TSqY0GDHJHF5kAwtJiUp0tAMUo5VKV+lsiQoKyEg5/GWx09+QW6EmJzZnshtz5nA
5i2atsXAWy6QlaAYOH/XOWsaoEohD7CTCIe5rUy77O/hSGmlBxQJtINbN9JIQdMp
LKJdZEpWqBv4KTAk61rTHLUikdEsPDqcPpG3tCttJX4xavaJTAjU5Rgi23ZCa4d0
9t+aGzpiUT6TwpZ03mIoB6jlNP2UrxDahQ/oFjUDqx7UK/A06pguYmNPQ+Gyu1hL
8obOI6RzMeeEJsWkIyrQ0Iqf8huD/ov2idCIebafnqVn9PNYqtSMebraQ05iis6g
/qwA6EW6VGDp5dpf/nV2wDs+UH0T1p1rSuHTH6eiO9LzHsTrw7y08qvGpcYjnmAS
QdTcE7OX3HDPKAgFWg9v0a0yA7ptMPbs5Z4Jp5Nfea+Hmpp1ku9xDdokZjuOZg8y
rQ/Z4AVdHjzWrvKASGSrq5I0MfNoTcTQ8558imEdUX7QvMLOs8lQk4itOh8GBOnl
Ped7svMbJrhiDvfsJ6Z6UqNPPO7kVUWJMf/XgEaEtk9YLyVzvnPyeWZDBGFFk/Jg
qXxOjwo0l2wetucVzE6GQ1aH4N3r1dsT0MIvFg7GNoNFhgW4j3vlFSyYv81YKO7i
Bt7GerlJSnymlg3LVZiKYPfxyMVxMIbInadA8ylITLM7iO9ujKNw31yPrwF7TBeT
t8gD9UWTU6sOOVXi12B7qCpF6b5ty3ghCbKoiYcpGNy4QvgV6Wk6QonkeuItMht3
av0nE/S49+509vqHgf+6fAEqsgZYeY25Jinrca+GS9SWUdjhZqfC7O8BpdsyGEQj
UeTMrvOfm/KwQEX6LBxBoreCgzrq66IKjSu4rcEp8sspJo2hxllt+Ad8GwPdgsQy
n+epzYIVQqD8EWBvnrstftdG8bYeLEG/ZY3cSpk1u9vpfLikN9HfQHyZBa2RE+e9
pKIbUXduUjkwc+CqU8eFeIXvbw6MyMITsa9D/VKX3wuJFK/PUrdR/kd5LBrpPlTU
fcYGsnpaKpIQ7RPOh4o89fR53ysdn0SW/Oy1/dHCrn9osS3rEfXMZH0xqndczGrG
hb2dBZwL7wZLinZkttkgrCk/G3qwiMx0HwMsYsRTwU/FQ3u65tppINpDR3q/wCHv
yWobHxXRY5wRmjcZTdqZEH3hr6NsURZgUW/Sljr5csZKnciXxqMfgRe15iXBlpJI
XNLCRCDa6ZqiNl0sb2XkEUHvIwWyG8f3SK0+CjTwigAMS3CdQ2IEifgJfdz32rTv
VCclj5G9F0sJ934audWvD68uRMN+w8K5WkTa2X3nzfMPBDpT5AK/RKNvwQiaibL1
5nJ/Zzbz5Ph5Gw8o0pRhLIMBHpldDqlDA6/LrzJfnLK3zBI4T9cDYN5Kw54DXTU9
IIZh3eJJrwRb6yRWk+XsjDWCy63HZJtB9TiyJQGQ0oaB0J1M+GmKBJhWuD2kGW3Y
VGFyMI2sOk+GmKllJGwQNoC2hQltbWCYwLurnAtpGMRzCfOB9jGuBMvV+4MUbKH1
27w72XQdjVtDUpQOgD2vtvvu+1ctia3kVtu7ndL15m31vU06c/EQLv2BSibjjH98
tu1+ElwBXIwqCc0Yd4DuMZ4m9wrDxjjevPwI+NdcJomKqLowwuUs0lT0lyeoHuYW
2XM0gFFu5ZR4vmAIhjlvWT9i3JvxqhOoa5NB/Q9DndeYmpvfZiKSVZfeUdp/kXyA
AIZHhkqXpl1+3SENudpQsrsrtJUgaZwMd/rypkoqeykIRKq+1m9FRZahhx979ZjX
PUVNgnmvG9Pcqlst9TWTXoQ/Tu49IujH/3bMlRFhu1JFccYvA1jY64mZCx2X1UGP
WNdixK0jhnpRSr3FObtvuFrMM5PN+ynR+Wwed3jBpBNYb4ctOiRq90m6YvuSK+cg
2nT4GI7L/uevL//nivlKnZN4ZzvYID90EQRJ7ChRZUmKhbN/VhUH3tFKsYa+J73f
2cwK2k1GmRleFG0x2ln7Dpla6OFvjz2UI1XTVhrcKKYv0nNU32YbQ5UMFsV2eR3D
TK454R2u4vyiDm0yzwRLWm63zU4LKBDMCLkE+HyWIHO82bUXuy4qb7bNi78+Mqb5
nuZNNhU06G3J2IKQCoQHYCPUN5vcTcxymguhhRJ3SaWuqBwqFL2mMtu2CEeYFkXQ
qPLHsNiDDOmAz/TEGQ6ljAHyam9oVDe47H71iAS9vRi7/XVQddObCJvpU1M4efII
/sBJBbndLmTJQtPeNmYl5zCGE4ZROdgz57D5ig9Cyv+t9mBhc2YXrr8W0/FOCdmr
iR5opSZWMCFwDUt6OxEzbPnN92vPI2UbYfqExC7YXU3vJnm1r5LRMJd9t4LuP27K
4tpVQ3Z5teieg4BQ6c8tavRsp7kh9TDbuEAJtCdkEjTkSSx3HLhDaR3MhwEnW9rF
JaCI2TlFZltQbfrJxJK5NtPiJ/0xjF3+wUHI7/0ufyN6w/vCx1+OuFwxyHqbX1Cf
7Pv8fiBHpOEiiotY9cW1vF/aAiV8bc4lCZvW6JwvoJKOKUWT6drEmcMnWe63M+V7
hXAYN3ObTdUEFVw+jOAqNsPkS9HblNadsi1rnJWHzBdP75ZxYCvHsj7N7GATX39b
veIMR7BSE78fB0+u9RliZ7pl8zQzdbr/9DwXXfCqEt9GIUBtyP01e7/MSw+ogocX
26uMT3MCRSXMeVJL86/PiNN09nMzvaVv53EyOZTvcfAiNX4Yw/swsEp/yKgYxtLH
bYFUbeLU2b8EfwDmAWAsv/SqIPkRpNlwnAekdLa8yXcwPxZp0e7BotQmoO/IH340
+NUqF6X2NQ/R2/fFNm1n/3qnQZIqHZ7jmhBm4YopA4clov3fG9mSrFuieu9pfUMY
z5Vwjzb0Op7SEvThkPF3IYo8J1oWG973kj07tylEq9sIpLXC1g6jr5ZUcypBHN9K
MlSOAEGbx4LQAMso6yQbqiWeBKjkcHv9Akvum/RvsySgp9dO97DZqZprqcTEo2cv
sQTQBUYGRigQlJv2+OT9CdTJhYhdq/EIHA/ijBKVmpXASeSRMbOIRZwYfB1iUnwK
fmNtf9d9tU9wFAt0ZTi0X65yREvwPoeMtvezm8g5gxlp9ZwuxUJF5Gw6s+RPA0M9
BdEvryPKCQ9iKRSeeGli3KT4oU6eMozCyLobekDGNyycu9LeVROtOOlSmZkq1cSp
8qE1P3fDuuVvghYr1YWL/PvzqAgtrC2/kHGMShexmwcNTvPLI3jfeGg2aWg5SUI3
H7DmHKi1H9TMD4a4c4EF+Whltxqg0rqiXhEweG5TIfWl1R8Ei271YMZWNAL0QpO+
Bv7s9+BV2uG14OAUajoUN3NoPJ/+R5Xa57fDzbVS3j734wabTLeVhO3SaLPwFyIr
cG4eZ9JeVYY79tfYl19xhT3RsQd8UtCSeEczln9PFn8mu84QH4I2ZRCbrxJi8mgB
lj5f2k52fui1NYsaZ6l+lCPkRrNtXk2DvAWKv09yoeMVsYKYfxe8JGdTcx4FCwHY
YirS9aYCsfmC1YQwtcYuAvLFv4jCwTaqC69zpkdsecdJwrghn3NJscm96SD0fFw0
xizE/7IGl9LYKML8ENVDDDPlItK0Yg2cxl5P9foiqXyWmSSF/SMxKaiM+L4dzJ/v
Rt0fQrM9D1FpfveTCJhOztt1cDJEfOmxfGI19BUsfj/32ta+9wSlmJ1YTcAlISUE
up4cb8Zd75KecFgOzuHRlp+av9UWYOa62Qjrn8nxwSD9l5sdTYWKmWI28M1lqt7I
BPNPeSM7aFuMmpl71GytC89pq/BOyBT1EPHevzemhoKBYQCP5xaPl3LZMLzjFV/P
0DztsAQsGFwUGfofpbIRNLluyEXHNRft1QvdrD/o4yjibD36cdAtkELCPJyByreN
zo1V3SpHrvYtUthQVYaQhM/qq3ot34PM6Q52TdGXpdHGWzLazKwM2MQ2zurmH6IZ
/9F0tDxWjndIxbxQNYhDLO7VUzj/AoFTHONHUWXChkhued/Kn63MFkGETQI5KeA1
y/spCxrD2QT4a6ay7c+HD+tpnINUHxUwosjCOvMoIC3pgr7IWonIzoEgenBAnkpN
lpBdKHk4uxjN0Jr+0qChlH5+MCA6PjTtoDyq3juPZf/Zd/VDvHj8/ZDuxfn1CMWp
I8/6pxLQlqbyxAEVUP+hCYeaW3fC9QN02YnVoUc2MLJwwLAzBYUss3KBQN33wnDn
7x84uwW/A155nuktgBpdp35SklkuZvNz1bEgvOw8L3VA7JqfQ8kPqGxv3sr7Gqhz
HVCLg25paMdjQ9xxWcqwyV0Ble/OUxtdJXohQWgwHHJmjt2OJ5FQI2AdKXwSTpoY
HeE4Xii+MmfoGBcIRAA3qDTU+UpbIZfNtRjyafPfdkGimRwMhTf2azNuYJhdQNmt
icYfkCyTeh80xzA7tF1h9SP7lw4uqWqbMJ9/gkrl6XYVuhek1+L9BxD+DyE4z+wZ
TzvmgPb5B5GkIMJD3jcu7p43c9H6kzodKf6C9bpLFe88342AJeubxucFSgegEI6j
sQVSG8vbuPArZa4RxY9MDqnUHM/bNnrLKgoH9QtSGL9VGR/594xu4QPFjyhqFv5c
ERSTRPib0aaY/b9GvnDO2HPGjwcOyhtQKLpgJBb8Daj8CbPJ8w/mA2mc51NSxKMo
kCorGiZEtM0b7z+dXI7J/t7r807ZFv0zFdAqgZBHJwqspR98QwJVR9aztBQrCY5u
IFn/6JLa6kNVfjWUcmYRqYbJ9SfyH2JLpWk7KhgmPYFRFdyq823qypwuxBmvUePJ
q/GfCKvNjkEQWJtkuv7m7yeXhts3PhbdMXy7fSfF4Tp7Lbi428YBiPjecw9q4wwt
XFlsJkxp2QfKTSApTo8JC2obQiPfioiwN4TgfcN6sw11CGj7Wu9TdCqezsMTVqYk
yTnjaf0kkzQVb9oLkBw6fcJYguCus4RAIsXm/2sGC3gAVaNLoXnFWT9n+8XCZGp0
V+cQOwy/OW9FG9LPOMnZKLf7udgE/sQeYQ0xgx5mmOQdxyV6A3o5KunkDOEHMnvz
DvfGvgmw5PEI1mXhzb05aTr+SX3tRrMLS/Q5kgI87yYWkYb9DHty/oojeCalQtFt
8dCUU2PCM1guJS1ElP/JjoaM2EoRF+jE4eok+tA5ew0gRtYqYQ2652M5d2FBxa4Q
5TbSPX3yflfLm63CLWrsDWgysXfiw7N/Oq530GivIrw3GimJn2EEYkrtK+pz0HHL
QrqfNjL5Zo3AFVwJXPqYQWVdS2JWTiOuLE3XjOLw/bLoE5lYEFhcWW2m2dJLMaF7
nSR6D4q3wYnJV8mLZLyob9i+U6kIeEW+scUky6718MXDPYmvB2HstM16EvmEuFuH
R4Jb5NQWEDaKIn/6bF9yOGeotsWYYFI6Y9qC0trVdfdALjr/2tDVASXYopPAtX/V
eVD3sy4rReOBcH49KZDp8JdRqzU+4NDO4Zf2UqYJcPyx6ZsXP594b+shI+WLz5At
jXfWPJiCD1gizttEpbKRzJCucUgDSYmMsvmKzxJ8I3/Zp0dZPv6G0rpj+HXjQ0eD
b0WFP1pTeL5M9YHJ8bD4ul/QT84XVYE+//uUA8sgXDZwt/0dw76wz4/lnr89bkgc
TYbk608ZRTbxRopry0FGc+DRi2wAFJ2e/YY3wKyaHYckTXxRNQXuakKCTiTOKMvT
/mWBPNHRZ361RaSW0oUGBSp1YXQo7Lz7qxfSnuZ6gm5RERxsVEN2BdrZbYLGxUJS
EYJLfLNhoWGyIweYtrQ5wpmhuWZ3DRklX6QlQQvCT5v+tSe6GM0gT9a5cwTM6RgE
OG9CPNPVVSFZSl6nqQBixkQsM/LnPNzpL0U7O4RI4ugCTaDqwg54yah1B8imACHl
3UtYJJs9NGLmRPHYNcHbaR5V6EdunKk/TbdjyvPRILh3UkN9P0moEA+Ji68qVPEQ
PGwjwdJH1qvJKaIbGj7YzU18W2BBpVyvgtH8VoW77/IF0u0KHA9HlRTTrYR7sfgV
eUuS8tCdqEh8EM8i4e2UrGg9nUMVlxNn4rLQfR4/XBZ9958xQN+Y9vf/LYn4gVgC
4kvsoZFhqG98SRLcs6ZRAuiuvO5z4jzEd8aUhsG1fyf/+tcO2YYIyVrj+uImLV4a
oc12ylPPREC9nxb/V+OOPy4btc1YvhQc3vVJfvJEOGGJpkTw12kq3+ElIMmbbSKv
9nAIWHRy/HGAviinZAQy2S/Yvn+c9Ypjm7w2CIVVkxUBtyIREo+IQZoscp2bfGv9
WbswUqzpJibaHgxP79hchdrfNWJ+Et2EM4D7O3inkCxAF9YaCaaWGzPoP+Kl0sf3
Vpf9mxTORqj/fSRieg19wPl37T6Hkgp+cKLt1vgeiFpvvu9qfCS/YwJtOxMofD+c
mOalNcG5nX1zY0rTlxVOojwRmHgyu9S3ojsuO8o6QWD1emeft6BVGQyJxEDYHR1U
OXXvamjWmknZTozS3w3LpfbIceNFSuTqX4ocioyf2L4n4aEzLgt3iFmaEgSK9TU4
4AQRpKoVpfhxM/yo+k0UYJm32VLVqEr3BBVxplGPmUSwk3kqyBMwicQhBm20qnwe
AYb2l1U4YP89KKPJm7cuQDGDR39nsRuCb+4etjc2Ck6wzhAIUHj1BbF3e6LTF8tZ
DQmSC2LHtrCtjJp1H1bN94GV6SaMEg2WuGEbPbwnc7e7UXrPG1xynl6Z4bhOtjcv
urtpqVExnUBUd3iSCNiCtxLv/8WqZ6qp2k+ywjQZQgELJtVeD+p7AwQmQV17cKdy
vlVCfxWs+Vi40LzNL4So3ZEjn6vt53QA130rsFOLP+R+hvAqK6rn829vYtOcu3nx
uusumOgqeGEHYq756F7uNomeMzkx/XcRbq0W2oQ6Td6yfESo9GzmlF+40CdNMvlh
sdXtTp++LOzYXFUYINz+MLJTToiz33ZV79HJF/7HWk4KFkENPyy1FYrn6tBS7A52
mhRSVlTv/SoGFJP0do5yU3fO+DYX2BuiqEWTGp+SY5kBVQfFA7htnkMFhDCvrmF9
ejedy+h1WhBB6IdNDC55L08siiF+4wUPCCyn1NMw0lLcUsTab/bYGuFqGU88VELB
cppQMGV5jwCsWsy+gvo2jMz98GkzqHVeARieWJlnolTxrSGv2FHvLZJPMsSqYquc
9ewfv5rZQlviINKSyDKlrPs9HUl4e2UnZONTn3hJef0wsI5yfRlHSpsI0CXDDEes
bBaznqiYKXnLZVVK0Gy7zgO2f/3l1FdltVlVWx9+ReJUGTMoZkEOX0DsoVBv1033
3qZveIkGF/YESfPy0u7VqlAKdUpNknJcg4Gp/VrEpvp8R8hrnpY8hQt55XM4v+pr
Gxeo15+IhY/JVkJDVmZimMP6WkFagCkaQKMZkvtKtYJltYjW9G82HZ3Unohtp+Hf
4/fo7JmFpvFcD2WRTXMokH627hI6gqdxrbVzcpSNgD6dN9vUgIIT28VEvdT6NHTe
GRXYImEw7KBZyWz4ZuKAKb2DDoTY1dUY/AJ4Yx3405rPFDzPzUxRohyd1ZCdmuA1
zJT02c6vw9fK6midha8fm9UEj5/HBKZCjlAZ8/Z8ks3VtA3cCmPhouqH/g0SW5hx
DZ7zpSIBVcO7OI5LokKLmmOajWnp9Nt9keLDIp4y8ZhNW08ehEawSeLOUQYn9QEl
miaMTAo/p2a81ngQ7XTAUlRwLkLgx3H3mokpgQZFID8sOlYcAHdxFSQMejN4L+L9
HeQDqLKg5gGfYRvxdGcfCmgbg/FEf0pao6BIDDkZp6K/lfz427xLxHQfjibbsMDV
0RsdGZ9GUkvzeWoHbImPDWRrJ7im0jqPBzrhRPNxXGnFjPs+wLn92OvPEsfe72jN
pA1VxY2gPbUrn5EtMX4N+Iwp2UPHgvO4wcvCPwI0B31adxf/9f9MEMiiWx8r0TC+
FsCyBKvSbCMJ5Y5U9yMp083BFHfX9/69KByFSRz0iJwt7sO+MepMZ0plSEmYe7Vy
Rjl4FacTR4q54Jw8C2Ulyljhapn4nmLHqgUlS96FJXyxbg4Gwi7gYQ7rpLpA3ZOb
qSB4jDlBATpBVlcbGeuiKCQ/PgfEidyv5a9NPaGYCHhv3Boeb3UwC0iLR08QEK33
ng0kKxjYVibDATmrhllP6u9i1AxKiYs0RFmkgrNTkw8fEzjBDPPbQiMAr61L5w+G
w6lpaaygBjuhQZJ6D4vpZnGYBnksMxKNy0ds2/r6arLI9NnaSzw2AhHwSS4DwrSK
G0lECzu/hvKy78dFyN8ucZd8zvI1hH1/JZJEZYCfboEFfEsL23H44RD1Xa8I7IyD
L9motEnpYEAX+lqaD9Mkok8kniTwnfKdFTf9m6VUcO0KYmbpdTVdIsdpNlnxHzHQ
hTgYW4qKE8pGMvFYtB/ukZLas5Q2STpruignPZ8ZhZQ2vKqjjkXmecYRVF9pXXtm
kaNbH+I21KJDAp2Knm6whhW4fgwXVafCQJzkkns+AIJC++0OAXAD0HTXQkCC29vI
mRQ7ZG+m6DkhG3Q/yGqUecdMkJM+73N5y7bNXubMXl4Q24/HotLwLXs4o0HN5my3
GsybA+W8U63YHRfoqpAUVl/a4j0rL8d9H6SMTEGL5sX8PT3yTxE99HCdNCK0h5Ua
JhPGKqWRNdaICRyW3fIlqhwSWjdjqfcL/z79F+KinDxlSwX9pod+uXvVozlGvn2e
V+Ye7VlD9a8cZUKrNmOa2BtG1afLCjt9TK2SclAneRgKnx0NzkMLaSED8LLDk4/b
yJKba2EldCfwY+IsPxmwU054cx0oUUX4Cez7f05C84ZJ9gK0Z6WHCMElESbQ4a5E
hSIWZ7v5a797dOr9uzieMfZQuByx5dpH9D4F+TJJ3lefgakgv5P05lBzcyZp58Uw
6KFXcSaOgGPmzO3C+ZQGfY1A4s3lTjTJ4ZE21SRExa+b3kwIGwXljaj+X42GT7PU
HryO7/ZX3zlUhCSQY/e60gvObBExR5U3o1o8d+OiITKfhp7kFJ59uHsXSUDXtRwC
MZKnl46G2zuJ4H5pUnsfCgIkVEh/GfQi5DEnxPSxjOqsjxkjXLBTu4VD6x2s6KKQ
jp4jxGYNw3zzOXBWye8pjhfxOudW9HsXD4bfUT2DlLjOoDZ/H/DOvgCYHufj2hD8
A2OSv9iLDX0Sr3Eo8Rr+f9mEwAT3Hlt3nXItDwzG+QmKLljFVmdlvqVCsMg4ZmBK
ehbeNLyS6Q25vwjH/v5EbC6fDf0Hppc+1JZk4Si4yDr5hlRmp0vtDkBpsPeqKpcw
cZy9BI65A6RJkDd58ZmfqjBWmA7Xn2Y0nb7jtUppPI4SgsSz7/3bg4t4T04pl7Cy
BCHvOyCZn6EfBcNcVylay3E+r2t1Ih0rU5QiXM8mor1+9PmdYuC5mFv5tSpZFC3W
ghKYQH0YamkfcczX1PDbpHxXUn4HCajt43JDanM2mFfwZCO60rR/33LOUob/HhbB
sKEbTRbB4L+zr+nll2wUmgsx451UX5aRHAd2hKNmQn63WDVreYgoydrbBu3wVV3F
sRGhHfy3XjScerKiWe4wvTHu+lq7gDn4WPGkKzOULaN08DvmOngQNgVl1q2Mff7p
B1L3cO0i9CdCpA3lH3dR6OkZu/ymMIloVFaWKQhIqyuv8YCV75isSZVwRvddUXBj
0Uzupbvv7kWsGQOZFHTUmnOPBHfHYpyiSK1UbA41EMOf5MJc5lYqexyXyniSTWwR
/Z+1ZM79uB0YLNIuKaDiut6TPdUKkxI0eOA3vq1teYLIFfWXqTQPGsEBbAnbe+Oj
KfOa12nBqvmcnGDP/Sfqu9tkFRlCEuNa+K4G7KlEaXpkHjoJjRMZNX9qnSyrcDCl
ea6ypdtTgnKkHgwe0PtO7gtqCT6W5CW11AMV9BA7KbN+mICGlgH1fKGQ2mdItXFV
++pIWOevXpYSmjo8cVrz8C6ts0VjJ6k1p53m73tlEjyB8brq6P92pSmlo38L+pKV
ZOfqehLLcFWlYD96qzfFePvsfrGoJzSNA3iTjs4ZFW/YPhfDL4nExgdEVp25nzi6
1QeBTxJT9+5rrEC6uoC9V1tJ4+hSBssMp6dLY0rBxjX/oSINoHnKHQ5KjIp3e0b5
0YTXb5+SII3/frHCESznsnuDLns43nGPrgF8fAFrqQGlV2YbQlFUOV9Ihdeo3Tbu
FHvCmsTOnCc4d4IVNPzXbwKtIOd7+0zRgTFEFE6IVxlVAYo+UEHtFb6yDVywME1A
NKaEi6HXYfytIuGdXyQfpci6uB7mNrsUlWB6wooKvg5u6W4IYky4Bs9t7Cia4THe
lneC2pis0ZCvM0StInizGemoGQMUpPMtdstI4bVgXZrLek3QCef3R39veI60bVwd
hugyutrfFiUsD4rK2g+14ED13anKymsgmT48wR4vh3HLYQ2ewqIM6tCRqB+jkG/j
oFLQJuCWqC3ZOJs8zJPz/MJfjp7i5MvT90Ps2Uj3ud6UyFa6Fu002yRpHG7g4U+g
Rs/Df+EVhPH1ON0fz/ayhszi7nvCdJz/DIXJrkXWDdR3W7jd2A5qtnbEk++1kUZz
nJg7pl8Ak99RRheS9aX9QbBfS4rv59UkDkFW6m0dr6jwrlHwbs7SLY3sOR9zuU3g
AhXIttkHwbSbpp8zuZ10trH16/u/cOWnldRhtPctG8u5ZsNUTk/wdBJO+PQMP+f1
zSpob/CRTJkhK2meH6FOlHGa5dif6WCc+lBGjm+mjj4voKqvKusUa3i4ka6QCDOS
kQA+vy/PiVpBktnzJ9qjmRHvf3JJrLigGVT9la+eH2FIlVmEhvmVef4UNZFrjv2f
V98a1D4Rot3oUy+KGZ6+YVGmypv0JA3vW8yiI1oXT3SLlsgaoAihyKmrAc7foouA
xedFU7fKCfun1De7JPRQWOGkTj/LOEaRvo0AfIrVj6jP8Tuke9mcrv7jW2Dgyajo
xpMtg25z6vPZFrytU/QlCMegH5qUXPof6g/IuI258w0tU45JsOTao/EmRWFW1Wby
2FyY0af7sd/f0diDAaHRLsUTGbkLMtIdh78HXUdRtSKHDEfA1MO01wEUnfEViiUR
0EAireY/wXDbk94d6mtL+fUbvSU1Mf3MMKeMQ3Pfz1l2QELUqq55weuChSqBB3Oq
fj3OOvGz9ICRwQPQrNq/coDl6hmrSRRvjJGpJ9dm5Pc6CW7uZlXIQIEHTFr+dc3H
twjrjcIN9x9MTIjzIV2IkAEyTcemgUcl5zqbrwqhJK42sYhG5EUfxclidiGtHA6B
rHVUa6OqR91wt0lWshkVcxhgnIEbOGcrB5RBJms4bGzYPvfqAswT0kmDOlHC7lDp
tv7Bt86vuX6B4MEVFlu115VLQ0czigYW9hv0LtG/sD9FcjqcZOj2cDhUSKT09ciB
wtxZySHkoiWJ9q9wQMCaYJteD+v2E/KSMoA5EXFpbimP421R6TcSgJw2uYeDoL0k
kmrjtMSqCZnxBbH6aqt2T1wQaHGuKyT9yeTjhWdSRfTT1pKZkRw6wO0bvAyCcucA
b0pCohMBj4rPl5uuL2fyVjS7qkXdH+lLxrhAMtRyUhxgA0o+kSr625JkLQ6RuTYL
oamiYzmj9eakGAmiwAboWN4c+36HvQUBTx23xlG0BPLlSLB22MAtUM44Mhz2AtVg
owZNLNwuOR10h/SAb0oQk9i+wkUw7bgrNkPolm0i+hmWK8ztB0V5fTJz8iBHoL6E
Atw1cojZxNbAyGDQ7AIpu21LDRppfOomeQ9tAOa3eOMLSa9GeghkleLDdMOwg2Vp
Uaq1t3mgAYQ5ziQ7hj+/EjysFGSRWKINoz2YqTk3JIoA95aCWmK6AFd/2MEGRKcx
V7je0hkue5ha1O/9PQBGYmGK4x3GYN9iwcSXdZ2zSR42F8OCsrBtFBL58LdaHUhx
ZZbqcXKOjfaBwugmanw+egzWjYEvOp+RitaEGvXHPS61Vq1P9nVfman/8fFpykN6
nssKQMVohRYZO5e6tVyr3xKYGdIoCBw77sEmQUmbpgaUtrVJ0BGqz4cnjrrD8hf5
bgi6u1275KxQQt5DFgrjXREzfdoYwnSmfxiq5sq4dog2CkVhvCyc+LKcCXM39DgN
7d8vwkJMA2ZnpbqhmP8bmFcRdt0dz65WgY59AWjO8iAAtYr+JRwEXrrWlh5Qj/kd
GPZmkGk4LuGrgbDZ3nwXafssDO1nmnYND2ZGDKrnNOVqW1xZCpwQ2aCWIAJotEMs
jei+aT8fygPNJPnW+5YL68EUhSWlMju5PXHfF5qbSzZFLIIA6XQDpLc9Dpij+yva
Y1atSolinRUUFD5gGazh7loOA57lucmcH6V9yMfystS8JBbhcXbZHpQc7s0GqSNJ
agyAqK//lIKebk9SmuYXJA==
`pragma protect end_protected
