// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:58 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sG034W4tV2oAwrIZbdvJa3dkeN+FUOQhTM2jd/ph229NeHFBIDpTr7xunB/Xb9/g
+LLJhFOOrxK8T51TBLewPXZp8MxWSoH7B0Qb7TmaElgE+DgqpTk18YDd0BAVcERZ
m5dnxEUauPGbTKp/WuQ0gdMp8XJf15jVYSYPVadk8b4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9184)
VBTEuLBizLjBY+RMu2bw+J2AobICYsh1gmDjcAXB7U+EgzeBYQdAi04+JYHJ5Zih
gIOxDjVosf2fpbcFXIFr4rVShA9RwZ0oqQujqGFHswW2kQd7WLbefOygc5gAEdoW
4QN0A6Hq2jC+OQx1z41pIIxPlkIwxPn/1ZCfiK1PD9BC+wJUu7UhuExLbeS29VaO
XtzLtK9LHSKPdc8Ma6HiM5pTgdNxvn32viiRauaa3cMtTr2rGMuYVAg9MYsE2j2R
2J6WJV6bB2zE0imD5VhXME4fV9aKK2LlWpxoHPR9fH+ECVJEIOur7LdwePawCLry
XeRIqPWQYoLLqdzEUd30cw5/tngZ5fVxCzeDMZ7KJQFH+cwh2uk85IYe55DWfwbq
PObcy3TEwARl3xTZUzJwUhdkJHRwi1N7WiTA/7/nNzhNiKa4nVoXf8AoGqz5UMZe
BsPX7og/ggQdujZQeRSlrQkI5/B/kttU8Of+xmoPu1o97GOtdBzcdq6KaZgzIHRI
97Ko9PAseISUAon0a5GbJqSwa5dnTmXW6fS8N5z5cQcDxyAEtPkShi4pz6DhG8PR
BKtIHD/bM2gM7xtgOHBwHoVVvJjDnbLkoqdIegnH9GBa8ULLkl4xVGoxPITxoQDk
elUiutvgOzbWsiv0Zwzs7PR+ftk6YDfsQ01D0ykFuBINbCAU4+Pg5CBSVszSHDmm
C8QXS8D+eBUQzuIvKtlaFPvZRjIcvdjEtQeGumt+mfp+jD0n5Takx5YFu4XzLLvf
Kw50xtuBlwO25mcZ6Q97iCf9zDWxFWMRseTZjbBe7/X/qUeme+8nNbfLkfr0/EE7
t24Dz4IDkrmB4Z9w2cbnXa8BO5o/NlbFDhCVmOvtTK0Imv8iBuvRaQVtRTO1WXDu
a3tjqhPTW/Urdvwb+6lKi3xtMHQlFdmrpM7YqlBRLEEpPOJEsNp7u/CNDxjZS5x1
CTobodUbKS7G2QehpN9W6dibfb0D5SVoERZQ+QhWiogd1PKjaquw9VnngNrX7vQx
PTGuh2RWI+kR2FGCI3cYjTZqtkEDIL1lE0t41f6DXG2yv1zUI8VAWkirJhtk0LM5
UXaTPZJFeZMlBV+gz7xks7TLLUkIx+487e2AXZ7jTeMnjIMr1AmkTP8aUAejh+W0
MUlsfPm6cRWSfjNQiB9h6uvy3huotVB6cg3ugp7+QnAMKKCiD+IVK+PMP1ZSNpJu
0W4KdlEpzq7qy5QpMldrD9CAIlbb4eAuCb8bhKYuwU2lrruHNDOGZOX6npu8pQhA
dsAfcZ+CvnC/fYEKGXYmMxg6csDZFe83bNmh0LRsjCEZwhV7hkdJw0iAukMIADZt
yhiRWWc2Lfjtu1eENl1hh/MXcR9IgANH463rElxiEBBeoC/Q8taUNqoI9ZhIScfc
lAHFh8/5lQt5DeQ/nJmhfPkBrEQDY0tOEUXGhS8fJJvSBv3quKgsUxrgx6bBpl2W
gxGOzQeS184WNFH9NDLUjZlWH5bcNccI7UfssW3NwhXjhq/0FyraDBMWyQzVO6DF
ZjQR/WLiPS1RIkfMo5eHTOddoepCJxZLEFsnWyjT0UF3DLSVNg1VyhdmuACnmQJY
rA9FUqb4y1sJ1oR1mcXGZZanYe2DLUf0S809MEjzA57jdAT8XJTaFtlqmGlR5Z0a
lgXbL7AOKE8wQ8WuwAp0PhxHpqR/vvZ4fOzSDSDq5bSPjRrYqzl/NZJPV6lOSt8l
l7cARpb4Pe8jUNjIHTBPQa0Sy1Sv8g4zAqygSoNTYBkcV/PBUUa2Bu6aVeZ+JTAn
FhDJXVMmTXfN6H7XrOZ6vj7E6hER44EGOnwZmMh9fYST2aZNuz5j/WsuobbxZimB
GzgOtg5K/DNWJjGPKV1gS6l+AozDfPvAQ3lsrRM3gwlZ2Jmh85lgna+48ofctLk2
UJyMouAKSc7noda7NHAzZNlQw6XAO2FZRQ3ouoaUkRx1Z22TKLWBo2bkeAftkQJU
UMOT3ureX0ZipunfKSGtRXJYS1B36eD5FaVqjdWfF4gImoS3gWERc7djWAJSNjRg
PXSQpK6fOs+vzaY92Mww/8bcjKM5t8oHT8G+pFVkj2Md4eQeifeVO3gS6g7MKAgq
wDczlFZKa5WjLikupIzlLQP1L9nEhxL8U+0hgBPPqNXdlFfXAX+m70CygiFU+Wn5
7s9wOd+4tnlNhAkyS7pNlbyrxxJ2+Hh0nqgH1WSOpWSa0rD7rf/kawv7G9BGeGe+
BxXsa9QDdJ8rjZruxepHWMKyGfExTve9WqpahfPiCFt4UTZAv36rUyVR7pbqSr1o
2k4N8UqSx/AVz3FX1uELUXY2iodMGZlwUeHj5/Cqufj/UpK9xCbXqvnTQ+8Lw6bV
WKDrOUwk52rnAzrVvlPUPuy7bUrH4nH3y2s3ZaIBejCWfMIyQDAwkbVbbvsAvm0w
sQ3smX5vGZuJGsZfheVVr9el9nyTxgUDqHENj/MZXPbjf5J2den/aNUUGXV4F8kg
dAiw2JxV8siHkhVWTQkc1b72STueMLi2pbETpptMcGKr+O3GCRLkkv3sf9EDMtt/
P2dyo5oCfgJzJxAcLyRYzyCbV4uMHp1jZfYM27EN9BrQ7PBcIpS3MA2RUBxeZ64U
wHCoKhKiIeCcS70zthDZWnvE8ImBWH0BTdwZ9HK4uZI37wVPL+mQf4ByOq6CLyRz
mb2S9PzBF/jiCKRFDk6cHplFHB7Ftigrqo92QOYzYbGASdGgeMQLt9qByRb49I3f
la3SoPwclKlsKR6f5i0IFxVwwZLGUh00dx220K6BisGlQgI8ks6VYlgxwYo9/zLT
/Foiw3jhpP+0e8G3f/5PKapkeuy189zq9nE17Ym12qdZxUxgF/6IxjwKfvEZNCz2
Wc0kuUtuxns92XcI36d8jp4Fu+d2dNXDs0GzIlVt49WhBHeKp0WjMnkir6Zb6O7F
QCHx6Uf/hI5xhpiGO/pvyedlrPF5YTHrz4bWzr5snx4ujiylwN9SACidCBqJ0QXd
ALBCPBSk71LREefE+orHX3wQl7C6tHNv2TeQPKt96TP07uJ9uD/n/BDHeQmUoKuR
dBPGJb52Xpq256Orro0TFtjz440LUy8UyyekFSAfdLuP5gyaA1Ad06edWDHrovma
7iOtHgE085wtie8R0q3ZrprZl/Uz2Pk0i+izVBs6fjrHc4iwMfQGQvVEvVL67b3/
yD2uHt/ID+PVr+PM6aCUUuPlANE01MtDZTwNzzUi1nKGEin7mJ6eDdSdeN27RJdv
QkSaSzlWy7+cx1JmALlFF4UQKv/RRalwV3yMHb0gFNl9voQoODU8Q/kiKdBmmzfk
w+ZVkWMsx18OveQOF8A7cRX1Ge/rNVG9bMymLmbZX2tp8wJWvFXb9+tMJ8FIDvCe
lBtbeUbLkgltwvHSeotCmkXUpjggvMEngAZ/iRaqE55EUo/j5RUb9iUGDWLWeM3Y
2a8a/1cU8JGwzNU1UgP3T55FaFBoBT36tReT/WAg2m3BvL4m+4L5tDKB3tl/fe/p
jHC3H/IhlFEgerlk+tEduRYkLW0wIqr+xUsVRz88MeFyLGcC1Iy3gy8fw6NH14nU
XmysDYuEPDrIojTIFe90RutOSMAuoz7KTh5JTZLr1fKmHjN9Ykkhvza72KpFuQfX
F3WE7f2/Bxaw/0kyj3vaPbkhs5kh2xKgqj59A7TATuMpBr/r5lw3Ek4lvC1ExR0e
elhMaHtRsq9+f3Wd10BSZEQgbK6iJ31HKPmvLWRjBKw6Dokr3F180W2aA9z+F0js
jmb+XO/4/ip1B5Y6O0YwBFBQxQSExy3GTYQk2UpaVLWvzy+ks1onQAgCI7tX/mtE
rt6SFnQKl5uOFoR6Zq3kB0VpQ2j+04FVT/bObRBprBLMnc251/9fr/Xm7BobBGsp
PULAIQZj7fNvXnK2KD1BO1Q093gTac/aVHYNKVuO/CSJdYNg13xR+QcdLbzSmZ6P
Gc/2RQtKU+cPJ6/zv+hDKM5UxFtPk4DKVcQW8oQCWJuBdZsyJUZR1IvDO5K4U3di
bPzy4TKjmWrZFKrICuN52Tu7FhQ1/3a9w3ZQn5vGTCyaXMhjkrhjwKjN3KeNxd0T
5QWQ6ZXzGUSgnbe4xU4c9JkXXTjRQDqNcMjBnyQgWQvnK/YUp6VcYkquEqug5edG
7puZ99DLzWRr9taJoDUqOe2tnaDBjaCSsSyuerwSybbfiFBO48/cxaw1eJhWBxpG
E/1YpUh9lFaJOYXwvr9YDYL957D98TSP3Rl3a3Un/qjt8dl293mmHI3Kv96kbDKv
UKVUR4ZfR3O83hPS6GhGNHROQMNqw/r8bg0L/nOcx0vEZ+DkoGrnEge8olsEcyM2
eRk7MzEy6eocwch+4qI59/uwzec+ZfWB4Sv/U/1Ew3T0ekwzeioEnInJZlA1kulL
BauLJnoT0fQXj6azmZmVETvGV7RT3TnOgOtNlaqrTqro6QB495TKuruoOWhDH/ZD
BSKfAw7EiKcrXwW8ZrfvITNn3T2fdpeN0l52zRK/VGGulMNbQ3U1+vs6ULrP+W+s
ETDdha2RwcXE1LbiFiT3+7+3/Jl/WCOLQQN3mo4j5m9rrmsW7LtQc/JOv1uqOmk+
2dkXu5LkWlyKmMKm/CLP6vdB9YL21q8jcchXR9XUvORY9BcSURcEOGzvT4w/Waun
rHEMZmOPRfJwGQQ879GmjcoFyvJgOvij+4FwWRCSHAOJpc/aIbHbceu1qOq6I6+H
PPEFx5e9YDVTqxGPXli6dp/tiObRrHjn1nX1K9uUPr7/M43eOcijOBaYil2W22tN
Vvv+BIeqn95mEXvf7fzSN2z5eveZiApcCaYjT+lD6eGisabXrwZ3fj2v17t7ohc5
5T42DiqZLyFAia7H1q4YgT8hJ1fd54k2M846EMHzAHsXhV6nLmK5CxQdSUdt2ekX
/xqEE4zZz6VRlx74vMq4aJEXXAmXu2sI5DV9mt8M3Uo35AAiURL6xCDPg2sCbFpI
ZBj8QaQA5Fgb1x7BuSDQelcRyAA2zAlVcr7FDv2MbD/JjW8is3pyAlwA4rb6sIaE
LbdgPAGO1ev/Wr/4so2jdvnEA+4a5uaArs7/+dRsvCJ8ho+ndb3z79WVnR3FyeeE
gm+XKySBCa4/SDVL7Ols8Rjx797HPFiFw9QOINXaQHTuIqlbGGSpmG53gaVtDL2d
soc5cx1nwKjzSGYTSDUSg0HiAZeu53SVnieAsALFfAAJZwCz5yfLSpFAGVnrGh0J
Oqv3X/fq61oFGAZvSJOZxphSXo1F6JKo3ajTVn4aHLQXqmZs6z7LIA37s9eyUmj7
3ha6TJpG/Dr7rHYPotqY2127LBZAJ/M8gNva1dA8V95IfOtiB+CqE4+qBORp3/jf
lFqFp5erwhL6wPDb52QWhyplBwaJx7CnW2lHLS/qxFcwdsy9ydNKVh1v5W2hB9/p
C3yxXlB7mwWoyymlym2dhDCjReFXRq4bq+d4hQMoBtuww/gzw6Y2m7sVDUSR6DA0
nUiq/tOt/NIosMa7xOtgeuv7P1BZF6+++jM1O3s7zZTWcmPr2XQIK/eWr+p4gfAr
92BZcijamyBCGnziP9pbqy0ALWPbN4qOpnQu+iDRHPRNBSFk/fAhVvjJzdK3TqJZ
hMvXPV59v2RBGhCNUe53EirPxz7mEfqOEuNjRg4Le6Hg0gb3Tn5duU81vEutWAqI
zX4XOPuVUcCRX9v6X7OjNJVpno1An9BdnnZjNSEi0yVfCF4GcT1twXt7r3rWhDxH
+AAT3AsQJcncbowFD/ZPC46dj5LVkLes91XNR5ur5tmIHCFlRyEQsMOZQm7AFDcq
C4Tyvw823uF8MeEjhmxd6I5oR3gt+gvat+IaCZkmyQfeSYPazIPBRjy1Di+oAd6o
g5NBwjosJUNVnHUoxrd/Q4TDc2VMmwyZDjJZfMUUm/4+5smuDEg+JkJfYpWVazuF
dDdeDV2iG/4QwJFRZKu7kdJac9J9v166Gjgo+JekDguRJxE4AhsCPaUkep27eDMj
tJk8tAGlhsj3GaMMP3r0gW+HgUkwEs7X3pA5N1xfKDaCGhi/tmL+xI5WL25mwRn7
qxyQJ4nM9pN3mEdbfwl03g+XUtY1KPNub9/RxspKMYPU5kqjwjdDhr87MfBfh1Hd
NTp3ONw7rCls8nsk/uCLB7zzBcRsBC7FMUmJ8aQkUEYS7MZDdPglm8JgrHP/+lgx
MkMwSQh5AViveUKqrUlhpCbkVhWr0svKPSGD4j6klNDs7SBcB2AZxH1rFC/bSSOi
4kq41t23TCD7Y4s+tC4C/a8raLxcJNE//MOdMBIOZuu0Tln0CMvHWqGW9URKycHN
s5iZmUtwvI5Mw4MbaPqlBzYJURsCGKu3VqdmiXtkKefMxn09bn5epl0uoXHgOeMl
E5f6eaPzvGewokdp55IBb/QNqrAFnn/jukZAwAQeQmzGbJ7RlaRx2QDkapSzEzaC
mjz+cZ3eIHK8kaHGP/C8BE/jS8QCMijt8VIxkagOzf08Yyn8wGIW5hGQx9HvitqB
V6qv51C1uUktrRPGgiHYGoL5nSwjCmGfpberylkQWBwp1awFuN6bFa5SBlrZmM1A
EGNoPviYrZBXFijDybn1U2i+p4RI7BjoINvWIbkmcmh2rmhx76OxA29Lrj1BAWz3
RXZP8VhBGBPNlnycIwI2PqQibrPaCdDNGpXTnHBCcAee8pUBw2FjgcSZglP5+3Tp
UHK62ybg+RzgYIt8kwHCnjLtwOzPK+gAyKbdXhh/nhs486WPy/TJjExsX0zwbDKd
pme7bJMWRYIRdXE5Q9YaLL/6v4zMFp4xfQgBg2Rdvl37pJF+JUuB/fm8sIb/bC1b
WwhYXK4ArWI/z6phyk63cuyhmFGbghcyMc8LRKgWigKAG7H4vGmMHevo3Nhd9MHd
riVITyptBgLYu7s7h2UlLNWLA37CtFHdIePd9W1fSR72+zWg5+Q68m8rAmUxQjBS
vYb0Z3VxMSKHAoScKsYbsE7jnohJVIUi+Uke5H9R1L7h8Mk8TmHLY0RAjhz09K9P
KA7JynUWKXlUxVlhd/AM1UZjKGYQZEjIOgN1EIjjaKG3emJknGO1DmiybbZn2rxN
B14W2NywQEi9jiMRHt/pEMHXK2lYaOEUjm7VzP9TLwDrqnIx+9r62RcvdykIj34/
inh3CFMhkh4XsRXPsUrMwTPd80WCCz3RODchHdiyOzVMmm0DY299pFqpCA/cjj3e
nFEsikbKp8SJIQWnHJOTtZH7xMepa964WFcfHJdlVUELt4g8alGutCx5UU2IE+o1
O/99L/JPSo5gxT9btVEz4cyv/pSSGlE0CHhv8nmk8Plt7oxHMoh3BLz0xhax8NZs
Ztwtxou772qxJXiPZE3JChVJ+C5iQ1O1Tul39HgPgAswISGdXpyLLcv0YD1Fwukh
rMapqP3C8BDpFDQEp3W1AbCgI4NszXfTx17HDAWBocDBEAxmRjVz1GtRwauZeD2t
L2lCoNwPAOMGGMRj0ShI3uhnJAmszz/a9VeIFIkh2ZlwWHj2kAwHdLdM0ndE/QiP
RiXXwd1alkFlLvJdWbei2toKLcYg7nsks7GL5RdyWKDHN8g5+gpxp3sDng17v9Ck
+E21npY/F7f34UccXDUoesL/C+Ggb2lLDuKHv/mntbu7sszsP0wLEvO8Q4Eotx+N
jxnx7WMzTymtj8rg5UpZWKV7dSkzO9lnS4l11Wm3i2RnBBxj2tIn4MKsKt0yg1W7
5A7yMOG3P2XzdYx3Z6AZRvvJ462pucsr35NhGRDUbaqJ3OVsuomqg9DXlk1s3f8t
XatJti7kfwqohzFYECTvR1cY5O+kNXvzCByJ+DUIRSff8jbriQd/hV8uWfBLrXR4
yPQDCIVIym5WirpTgdsSuPGifxCjrhYzAi9K1s8a1NEnCPKK+sKKfwFgCaBsNzc1
ConSu656UYA+td81p56ubzDStdDMBfUx+sjdJ7wslbOZoMUZJE+Wtda1t/am3v0o
pGDH0Te5iL32fSRrH1KoifhhCtyz/z7KFnxWPgFOcuHHqXZEZqtUWLszyBRTiXyw
Srkepl0YSuGQdjKu8BYwSg8Eq3zB+3YkyvrZSqauBD3QYYV4h/UTq3SyEV5JWFx3
djOWwnq+y8g2AG0ddzIpwuAFXKXq7jYZOq2pPMBWF4SqwQrx1aayPfm14LbBMTHb
TvhlBN75tBRisXKuH0SiLeRdah34HPp7jn4rT5A6QvAlztjgxwEmTdmgVatYyPw8
wCj86S34mkrAK1z4QbFJxmFmpqaJoljxatMXCzlyEuEwoOj4leAp4K1zl7MUogs8
6aeWaTXfC7Seyh7bw6ybtjh2hu0YIi4tg9m4C43EyQjno/exLSuS6RzX7kCO8nT+
0/z2efjLiPu5LXICVQW/lE5r5wrFRQKeV9tzX4kPyKE7iSd3h1r5+164NIocGvVK
vEI8xTxXMlGJrXPbeuoJecNaw3t2oYtN5qEebQJWZb4QmgQD0JyLrQPMJImwq9Hj
OO4NaVmrpCm4fVR2TyH1s64cNeL0aYnKeac9NZOrVY6rvKiShXMvrvnlGJ4lC58g
EslEXlF/sKyPcgtBWcqIrDeWWei3DHJyo9Kz/StfE6P46QhaTeLIxKj7JNBBLHS2
6QseAis2FRHgI5e8f0ch7h5vcbxoRu9V58NFo8lTSVGd14XM+cbLEHpE3lDbOqUu
Pi9k9xbfEi+u3GrbUHruORyI+KYGqdlu1GXwbu2Kb/PNOjtrFRe4qrNIufOvRTiN
JNUk29cdolXvM4OceuCzcX6Kmoa2aG/3x4nGgjuUHMVjuhoI1tYulcTYGmmmklNW
CFCm9UmW8x/dF6IpSW9l80yg6Q26EeDr7gKhjaVGUGBdYBFQmdCWmhB4ygPvT3yp
J8YhtlECAeMHLjHwi/E1Fi8+NP6tUE/kDsNshTcbGHLAV31TAEdy4AaUq52/P8VE
P2zmI0VNdq08C8lWxOTFquRX52ph88657VwHnulwtq5q4XdDD0lNDToqzB11zgTa
C2M0XHcPLDl/XUJxvSJMiAjXxNfjx21IHsrD0uVYGhyaewbxOZUohWGpA0U7fYOI
0ao8IMpoY8OqY2Byq12k07KTU79z3+2BjnMFyXZWwH42Wax2j8aAjsDGXZYAja5q
JmAZWaGmJLLFydCvaQT5yxhxpNmVMGzBgcnfEQG+lFRUk6QsWkK/RUDywwy/V5Xh
o4edNADrnZukZG/M9ylSBXQX5w+HwhnfsO46Ttcy1GDRHalO3zkL1NJDBZSjgp+t
qrXBg6h/Z0vbx6roAxCc7yFSTIGx4JPXDRBA7szv+ZRmZw3aK8tX0YrMV37uz+DL
iUZNwlgA45xKjj6CRNGVjI0VoyB8nbH9PSdQcU1ig6IaKzSkCJ2ZY3nraw2Zm5w+
iO2fbczi7ncjahWgo4uNIpZJ2N627t4RfNG3G+id5jjU13NeVL4nH3IB1MyWVs3/
zQw7Gb5qK1zYw6qE30PiVBv/SiJwxqnBcMCqHQNzFBisUUvxQaaopboycGfRZG9c
vGRN93mvG359+Y1znlkneODcrMuyo6r1Ck74K3xQLcgF9Ldx081rINmAtfcL2iFA
efUFx3bD4Kyoj0FU7hkBysqvMr6TKjW9joxQbjnA1l0y4dIzk50QCcPfJNFdGhc1
mDxc8iGDtEJ3r9vaDEDYHfYUnx2g8Qa4opQPLVsvX4CgTcMg/Nha0gVD2JOfk/QJ
/97LRbWV/qKBHvwTog4MNhG2TKYdGrWZl/mgAz/DxpwV2xlh+PxTzG4OSErIxKXd
KE+bxxrA/x1TElYTJNnn7BRCJJP/rmIt9hDUP5SwObJLe0AzR0H9qIZgd4IDa12Y
tzYEWkk+VqagUZhY5JiB6NMILgU0jLwswlVdA0yAmEh2NPbojY183ABLaR4Gqf3O
V1VGPnfYlmKtHETrvpn+xX/u57M0IyOBtlUGQNFLXCmOceV+lwOvLi28wGMsG71p
95gOA2R83BkEBpiGJ5ltA+zaQuWdRUlOv4pfl7YZMvw96x3HXTb8TYR6LrThza7V
WvHe5nW62j4/RXvqzp0txN/hpenoQmzw7+oN3fWyQUn9fnwkt4W4PB0VYQbdHbfo
WwZ7KJItUb93LIjAqCHQRrsIJmiljuJjfbEOGOtUXu0Dt4g6hsq5HGEA6hLorx8x
Wabc5sYKsfwlAc4FvNJsUK3uhEpxMiCRQJiy+wI1+RMHasiV7i+oKQVInho1Y/vP
l+SgdtClKaYPI/cWmUA78QYTox6HunnYOKvRdBoBdJTuSFmItsHgi1r/yJjt65pY
kInBqhscrLLlKMWpexNrkMZuuRDVhEDhw355DRjIegsi2uP7SPah0PEWMdDP4NbP
TBGsrfxKyochYYBtRT4nklmfHGsfQKJ7alYjVffGePFF30x0uQtN20IQfpY022Fp
tz9HW4vqR1cnheaokZRDugJrCa/ZAOLfdlNvxncia5/AIfobp6uMxNYXdKn3DPC+
+uF4Zd3I/k14xGGHPmYTu2522cE1XPZ0tJYhTxUtK7YktBHYqo1Jzdo13rWLr+/F
huaIbk840pJuqiAaoxEDjRBWJOkT/s5boNVF6zL4VEwsapgGYVVmBZTPgz57ExSB
R9Bs+6otx/dzPE4JsQ9TBpoX46qRGbruNhHlVzXI8YVPXfpFEwzDbtcgKrS1/HpB
1KSa/OyXOqh1b6dyUHrKrkeVEg3TPbhUvwpG4IATnTdFDPiByLuev5HUutezrtNI
iD/B6vugNT1ssDenrGbn0mw97g+ZMtJRnM0n6hkY/H0yXrd8xLh48Pc6My/A3HrT
evIohhkNiMD9tbuS7VojHIclcELep2gSQJORfCHQg3MhfrYLlG3pGoYT4y5Jfd7N
Ue3GlpGXNmmAnutIWlOv9qbyNUcLq0nlEvau/okBicJEjyspeaA4CEPn3vU6awG+
kuEvtw5TnEqwoJvGFVcMxis7uM5WQfeNzkLxTcAHbRo67m1Xw/Tfpk9s5jTJavGQ
LeccTGk8GLqFV+e/ToaecxP5r/r1nVJJOyCQ0kpwOzYWoHWyDpwx0BgN14b8JRHr
Jq3khuICSpMgon1ELrctNU4NMZ5dP3WG08938oJHgnX4xA1rUmGe2EDjE9p9AKRs
jEojoDqjD1v+6e1rwBW0Rt03ZoEaIL2geb7JztBvki4QyLc6PQeJd+5paFg3pQLb
6FNnru2+xSUOZrL8elqoLRE9BjcnA2CQHKJ3K4Rg5Yuv/NFdbx/ELQeL1luM7bl3
MtKizM32AoRkQS/ZiEmb3CGeWIEIMYPYwuVUbUFB31d9kSF5IaeJ76Z5iyvRuvJL
EWdELs15ZmAzHI/QpsAa2952Lyq0ntOn47yUWrnmjMXejWPCX3tnAt/j4AaAABux
zSOmC4mEG9qX1OfmBLBqIXOIXgffaAbR8ZZsrv1L/byCjLfXLWBk+og8cgsrdg38
j1Svd7yFGLr5dZkR6OPDR2mjmQpgnJ0UywxE2UyXxHMzwbsYUaSt7/ZYoKAxNB0b
gZggRvIFs4R6VwrRbIASti3lmSw2SyjVDId5N03wKHfefnJEBWwONJaoPw63INoK
ngeDJ7ESoplA5KW2nlUsXLwGT2XUh5FELNqR0V12nkK2sWHEMLj+R6FALq8JpgT/
RoDvj1QWeXA/G9tkiuvrdOkgdY1ZNHHyEc+tM2aE+vJV8ONheG9W05qsiVKOGm62
/IRBeEQkNfwMMWfnfOvrnYMGWEiyVtR1/IS5gcjnpjduwjPVS30PhAFscNncnT6x
XmxkhXWgGBNq40YqhqlZzgpdYy4kyUOCed2ymEyubxJq9JiUkBY/G7GCoqKIKfta
rCbdHYlALOD7c7L6aTtRDNGlA/aTXV5f90oLYlTl4/xUEtFgYkgNo2zIiGORtGfv
Px4WCqc1T8y0VxmHwikoOubTeoaQQSoccaU7zjo8HwcmrbKt+VEHfD/CY8eHAscW
kMm2uqemYqWRtOy7TSioYD/IRiVmTzPZRYY/aeU/PttWCsP73ieA/7objztSo85O
4SBv5Ra9POYY1eT9mquwfi6tUe8PMRhfOge9FNDxFR6AHRbm2kox7O3T/eR2ZD8C
mgCmChbSD8QGX6it3Ub5EuR88KMRcVr2erA9zZ0zarItcz5MTD2DlPdeD3YJ2aSe
ja4uBmoYF/rW7Ue2UXjmCFDPu/Kd5CsYhYdE2tIXesXFjid2Be2tJvm8kUKAL0k7
7YXQDZtNtIYaGuofcmtccg==
`pragma protect end_protected
