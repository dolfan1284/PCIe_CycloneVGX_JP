// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:04 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ToDzI++6Z1u8bihk2L4+kGGm5h9TXmxEfAhOCkB2sBDrrRXebPzF2cRifGtrj5lv
CujDiWgJ8YAWmRoA/fiMVd2soPpAMmctUtzTHqghPKJTUoaN+VxH9pljrKK7/XWZ
23IsOlj3o7U9CRgfboSfWSV6jy+JTv/roD5HoGkgUtM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
aaD+bVsbuRJ+YYI6a8JY3596Tr6HLkfVlBMCoz25NEzziB1fKjgIyPIQa0xupfJL
hAAbFbv45AhWTAX23OH5p49vL0jsubap1oxK+KdAGrsLhFBktghnWaze+fXyXHW7
GIxc6bXHVlZwWN820SokmQ1XaYDpKa4wpLC7lILHrmSrxeDWajmvr72Ui7hL3jr4
e6RBOv49pUgXHOBNVddvOp/N8nWZ+71booi3lRR3IOaawBNCCyGxPHDIz1DKT79M
c9k97IcvcAM3rAmgG+8vUyM3jVWeEMVOADbLnkglndDNDzobYt2athfMR3o+9iWG
dUi7qnFy7qhcsWo9V9T6+n9tcG+Bawa+Z+mub5KkXGyLtlLS8aWtMmr0VebyI8xv
A/UZJuJyITRHIwhiGaLvnwKPLG62enFd6mSNFrl1XoNQfP7jJ2z/3PusiY9Szlzu
Tvtw8ldnbuOQVmRAub4S2ArQVSlqPjPmHWJwRPGmR26aS1NbVgBJYIFVaTqja+kk
5WAEXzU9p1hiXCaPwuzCwfEKy90blf9gjxJIhgPXrq6854JRpkw137QvC5sB2ZD+
/G6Snq3UI/+ElnjOqGMbMzJbPEM6hVzBtS0wH8Kvv4zjFMHpqjkcvATgXInrl5KX
v/tnv9QLdHIhbgOTIQRpSnVozxVMssL617rfddKbaYhHLgQNWYdXg8UF3aW4ZCr0
+INLCo5haS4NDR4U3z1ertn6YGKbfFGUaF9ifMUurhGiXDxReddgLTKaQ5mOCv7t
pUaDHjwTOaXFSQ7RNL1T0Fi5t+OeJY66dTA8Qnl0myUb5754yAIyRMoFDYr3E79f
qhIOgEDf/6+PQxLA99NwQqTpP/izKEO8PZyTuvuoLa4SjXEaOwG3kbYXaorexDJm
FkQqS5M0ja+s1m5dOv6m96NPVS0b5WUe+6fju4i0P7ucIqdQ8XUqjj6jb04O5iGr
flWuhrPqE5MgQgbdrdZsbCdeV7qjPIxv3eS7veeL+dYhqaUDNUJUdtm1JDMXU+Ar
y2+ltOOXoLKNCYY9rji0aKZtxeVJnAjc+E30bD6Wkt/N7WDs5D3RwhJy3DeIUZ5F
xH4zeY2p82x/Axme/vXgSMPj5hansvk8oPsCBdU/0c3LRy0i4GELti47h9DEf0mz
Y9wQbge2eILr9ukvO988Ccf3DOf73g+xOu7kKGzAxcrPfGSPW57EtMQe/9NvPjin
iv5pW1NVn0B+awyYuvQH58pPbiAMRLDYuaRA9dFEkAcqr8O8n3MX0rUo0nVYDV6L
OqZgvBLO8/jJXw5tbBrTef39Jd1D9WxEIpCYM05nySrY2GuvCwoSilPCbn+TeinG
YWbt7zD/Oe4QxQbGDv++mWa2GROE2/Y05D7n658qMq/IIEs5k1g1OFv3rO49AcSU
dDDKRrJd6zAUppPV3elnMffDQxIhDY/t1vrDhMdeXHRwL4N/d+IrEsKeNHcQCBfH
fCl7opjg9fV3RgI1ehXn6HnT7+wSTmYDw2jmHDcXuwALETJeBKVVedpmGY7rDQkC
t+sQinYzg7oZQhukun+8MyHDHFcSACHw6uLzJRW25J1Z8XgcZtpOV7QYYC07BBgV
lmRX0pOqD2gKjMzDm1k696/6XkJVsB138jzp7Cyjk/u8lVSy7bWGjypzF++4IsDA
u6UWTPzJFElt8Gjh235N9CZZjUywDqmqjn+c9ysz/GiJu3epEEjeR9+Rr4fm1QIn
+5anJon5ZbWq7yYmyJ7EcMgYJxrsKz1SnXuqLhhQidDOVBKgY8sxt5FCpZGmn+h2
3eZ3L8WX69r6/t0Utx6Nlr3460XkMCem9oYVXsoyVmaoDKV2J2T3WTUcd9PQtPK1
OnYoQC6fMduGsokWtJf0wWgMAKCtR5cgvpfrJqBFsUHpubesjQmtDnw0Mvakq42Z
igMgluLACqAJGyKSc4fklFNCr14a2J18ltDl5R/OTvgZKecXx/CqU6OvVYzsYLnd
ppBR3aYGehAe1YLgsJP4n/Cb+YXuoQZF042iExSsZmImYXvzlnz2ZWFk34TTU4HI
Jz1O1wnsjoPjAY/BxmBxtVRmV9iGm+e8KjR52T3+UKQYT5F2vXzSwfHpZojaxzMO
2eht3ujEjdegxdaejgm5fFm9zcpb+zFq+nXSCeDJXyAKlh/Is0424n/d56y9l9aP
ikzeQ0gk+EQNHbBQOXBy5aekyb+x+0mekzfr8tesHAM5fHIc24yVkyIj3V31oLba
0lXjKYZgWeW+Fz9Hp45aib6pYBDjvrb1xxtXu9Gw1q+Dm1vbYCSpOn9oR7JSFYCi
t0or6I8CpggMJ8xHobJrZD5sfqqCOExh/UM5LTNX9VJP/BZmd/Osf2MJ7IQHj3Gw
rSOWGRJ6l3Xm6ky88poLhOuc+NilDXs4YXvQM5fSAz0B2a/el1NAoEXYGsME0ZW2
f1L1XMUfigdctsqw1QunTjvSDRQhQUrNAv+YifkPG7pEhH2qkw+4hm2OfAf9KCgs
f7gQ0a/f66+HJf5ax815mCSpgSwq2urfZYo7BNnzoTAPCAXps/j5XYWG9uq/5WkE
xOo8O6163LJ0Q8t5kHY/HpJG5duv9nC5/8sfpmbEIBlAdx2ZqsDhNrtHMWAbQ46/
SFPy+zj738xHoFBm+1HTykxL24qEN2JkMzI7YncJbh5Q2DN2/BZ2uEIrC7O5i//E
ZJNTf3kjt4dg3OOfTqe82iEIsaeLtrVjGx1F1AvI9JAoPADypn26fc/ZFpQYj4xM
lYHQilq/fy+pEzAfnHL/7iuD93k3+3pUxBotmGtco203ARKiaEbDvx9z136QvN6P
xNHuU0J6TpdMhNi4XfzJs1WTd71HUiyQ1VRPS6vRpSxYGj+nSzwWQ0z60Arnq0bB
s8PC8Uklbx9K0Xh45TVQfA7ECbLYneni22cnTWf0edaue8fymOphvgutE9i5ft02
Uk+Li8YRPUhPvgGAkYfffhO0BJe8FIklrG/C70y/sDrRsNatZvlyNGJmYnjP23Rx
yO/JXKeCEF2UCeLDEXEERwOBDZBn1C+0xRwfK+7uWVttJpH03z3493obsfUTQowY
mM8sZQoVDaYT5lpUNtmUF6beuS1arOT+HXRjfcCk9iHgxoURQGgwfHOdhP8lFScM
GkqFeXq19PalKA85LFk+A86znF+3sn9MI6l4mYQjxUq17dTvksjzF54xYvOyLQ+2
ppkVcCtbzh2CnMTPkCUDbOaUWkJSVZYXVctDOlWSB2EoCCBYHiLbGH6/u7VkbV2v
JOVemFX+K0j+U6UfLa6uUXaNJ+FvXmQ2aY8UO3I4MLeyOwiGKcJL9JJY42vh1shD
RHzrO2JMDshy160TLyUu4MyVFITENfTRNiHDG7mPhahaBzSLwaVpfnbSWX0Q2Xb9
r2D69P/cd20oq/FlTJ1R5JPJNacsqz5yuK7ORMAWL06+l9VX+g6jL28KqIX/c6Za
icNS/stsnSIepA63DAlZo7K35aJ3ncfWjE2+Ruq3/hxrGBj128pqP2NSUPlQOrKp
58SpCaZFMyp/XxYOnvB6q2qwwt5u8j7tql/wyoMPyM3ogrkVpnRH2MHouJfQT0ZE
XSUDvGPFD1GH6EtZSI7Oi1mEwTmo0fE92jCSXR7GK3Fbxk/2B6GVEcKv15a3PXEe
Hmt7EZ+KNy1J3J70OrEemYRqbdgkzyJGdWjKyfyCkrQAugGQ0jhW9x0nqz2aDW9i
jylfeEjq5gaQCUOO50OhVMwcfcIsEIPE7pdX9Zzg31GXi6FxR6QjdzbnuLbaIzMl
PvKPaK3rD94ANY9w7I8RK7O5HHHeox0zFixm1ygQgs6yH5GF89PWZjFuiREcpLDR
C96lt6Cmu2MGmDaOBmaF1ZEh7HQAyKzv/k2Mwuti7PvWxmEKs4AaSoWA3I5H+608
emE8O62CQVXGV3H3F9Nanc1kZae+sxtLON46TU0wG6Kv/tDCd2nR8yXjcb9+eFxI
4JhlYK8+yOUkkU1ROApE8gypvNALr9uXyGT+k87f27uf/V8gDclescU661vc2+Hi
kZ+zvZlap0VZ3PICR874xBXqaxoEZeDmrQZLh3M47nPFZwAlHoo8PmTqlDQIl8QC
ZodPpGkTnOfswX9wgW/RXDQAZMGUfxswRs1cvbp/OOEMvmCL53dx87QMXDqgXSPp
KdkqLN00jadjRdL1RnsQB53BtnmUsSa7ZzEIxUeQSS2MYYhLe6DxLqBfuNkjYuWe
GT8M3ZiFjPI//vL3nHq9LSIXrG/S/nkS3D2YoCXifflqVZfOyAT301GZn3K0+cTO
cOpdyquIYTB8cOYRbVI36s1PCCwiiNNQszQ7Ct/tyPYiL+aKBtpgghmuRCHDFre4
M+CZl6yu/oSGn4tX8G3itvsFuIl1KHas7GL3av6Go7JBvgf2we10C/ikTf7LE+qw
S16HUBOKY9xPkVCwtyw5B1lJCi53e7X1xYae/N9KpSg0VbDkcEypJSC05jqVBhlg
Zz0CH6+G9toObBupm5m2LXROoto3uGYKgsDZeBRFhSa3bd//b/0P3mVe3/TbVzu8
GZVb8vZgG46k16SQsGpdd3q82ZiNRl8YVWHnlr7sHsw1SpqgiitbrRbX08sDEXbC
4NnZDMHFHxSx3vSiaSSJ43xeqPfr7eurMT4L+JaeqDOe2VnScYnmJyKDqJbLvPm4
26g55W4dpeDPyZxn3ppX9B+/gjl6Ov6BVYNJalshl1QXDvHP29d4kI80b/z8Xh1n
xYRjEJQJPsqHnnPH+aVLdIUrQb03HNlYRv86WQjkUPrTWIyLtxCa4+vAwJ1EXaC1
5MQa+ALPOkbBYhlu+aUUGmSvdA4GIw7JCYP67MdaqHtfxseEIIu3vClZuPd9VXf/
1vmK2+zJceTJglcdhyp0EOmSEZEXZpjH94MsBo0JQVyj3TZrlUlGkgR90AQFM/t0
ClV6JItvsL6EKQuKIem6a4Pr9hWwsXSPFFj0+TIistyNn6qJBKJkfq32WCh75M/3
G2qNWqzwZhGyjbtf5MKKKg+fOobYFQooGggdQnveGAE9gHcYah5xnwW6yGGk4pxh
8JVGG6uM1mpTodgvAKv9pHiA4b4PJgYhQPLRsPGoD2MMWRp8oGN82UQJmlbVAfIr
/BX1Cf8t1m4yJ713bY3qprD/drB3xw1bbemA27OE1S/uKW746cUST/c4QiN2QXPA
kvbo+2hiK296DwgVf77hSybgYlf6XrLlQLW0gz1CZvoMrHi2nZrluXQ7nfvH0MLS
Se0YDNST1xuOek+TUTfrvAqSaAOhha+BSIfWPYZ54FBi8PHU75PzS3PImCbJbwsH
tXsMtHAfPgmVfJAwfhOSg/O2e8njgf+UVXncMyYdOmfkV0j0/2IpfriVAovFCYaw
gUkIzJT/BhU0644PnU835VhlrRy3vtbp151S489gB694sqmncsg53ApCNxLPuneW
j4STYs84gvdaPCD9xtYSxRHNFb1bAZl+V4t4LJws1/1K6537UPQm4o7bMtbyaT0K
vjoPb6sAMaaPVdhvX5rN/y+vgm3fQAcjKw3ji+03AEzB02b5aqOId4uy82KPcJc6
MYsK9kXMoy/BVnlTN5ZKmvVt2chcCkykuUt/jcU/mQgS7C5/brFh1TgCEc7sC6eS
RekUHPF/Y2pVdvnZZeLs1qXxpkaBa6wb6cWQz7OHOF72Tb1+b03uYvVdThscUGvR
wCLKrY0/OCr1TVtXta0A2CiauLlSDXWrRGbcRnDjWjtB+LiL2DJ7iBodQW/bDeKn
0neLWr0VJzEwqnGmrgeyBFSun8tt0lRXSbJlLPn6rSzot8xajHnzQgbBX7CkMJXX
NhmdR99oXzmt9THIMpCH/SGARMGjbKFpzRLfZPklB/HnBMGhUvf5MLBUnfYvvTvt
Ps/Y1z5hEjrKn0B46FiWqstsh/lscGpl+cIzrpzp20DrRrXITkXb37r5TS13dtfC
Mu03Wne+tq5KdIrht0DJr2Nn2kslPnLFHKLc4xqeBdD0FADCwomvfRgqEluXLDNO
WFYMWdeQ4TuJObVNOeZsq4bNt58cf0F1IRkCG3rOjjkWR7y5YmbN9QVb+X9kvPW1
GJwjVWK2NT5zhgkEIsqQECZJQzQMXgg55OCGH5kLPj7XdQVVtEp2xlV+CchPLnzM
dPEy7UXfMBMgotn065tRv5dazn9AUVU0PlyKFZ/QoHW952iBsAbKnEwOfvm8ItZh
X2LWxuBS/Sg61W+RibVPZdCBrmGCJpZ3KbI9NZn+gOxhYb1sZE+Lhjh+kDZSIib+
V0R6Iei2ydm4oKnAySM4YE99+ref29gGFN5+8SbJvaMypuedeHKUNBzDc3BzXGM0
ivykevpxVXuOrH1ePNS7RQP11IdkNiDQt44o938JkS3nC/CoRx6M9hN1aXYKkXph
NTRO3M+DqgAErSufb4g/HDgjdEKckmikDN7rAFktOBEQKQkpPYXXlXUar8m76b6r
hx2OepUsjvpDNSvZS29v90srWTPtjvYcGs5UqW4kXXiUpks76xbbzllThkjdg2yC
XgSjrCL0xMvi3UPqOHHgiS6ODmOpsuFHw066ByrzNCAA88CPmMTFC1wiuUw2a1bM
DblXEMZvCwjnOgZWE+AMhPPsBjjdM2s8PD5Z0r7TW7Z88pBPZuWPmiZqgnN+qMqi
oRjyBauJlYi/g+hC43vOXNo5sPjymJyos46K9UR2a3IU8wn0vyjEE4plJIsQWP6I
34Lr+iNaBQXmlF9pCZvHwUc1kw67NiGdy4hwglEhAezoCF2TATUgcwxJvnZimXoU
jAC1XrAdPC3zWBPwp+CJ1LkxZmlw5/iPtYwBbCZgHm44k4QkZ6vuDtAqigVLSM6J
VIoSXZGjrN9XT042a3rl6kA8tYC80iZHd6ANwDllF4jOGyADRq3jINduM2Agbv/H
PJ9OKp2WD+UUVBUNGHZsEcXjO5/2ni9nr82oDmqdl9UQ80uS4+sXBUpu7OMT0cIi
Agfa5/qA5CA49+AUav0YId5HmqPuEWlsKL04rmeqLGVJ76YvYEue9LIDdRD8OI1S
4oOUjXEp+0jQA1XL1X92nfmWWpWKxoL1Xaf/mAdkktlz+H8G61mqJwPcNblTGh5v
o1G/4zZHTSKows7Fbys4JHXSuEyFz+o8FraFdU5pY0bu9LS/dpZibP70NbbFdhCu
f9trOhLFx8vJtcAXMhtysgBuh3gdAwsgTmiFh14UGcVrla0pYDLXd+jvFy69o/py
KoKtw7yTpiTH4iGs4rd8MUqfOaQdjbpQY8SfLzXjxEIofeRXdUYgB6CH+uT/xFvp
FBffPiycwjNAC1X2utHUoHyICbbD4WPwuf8SL/MnGp9Mdv8/FUWZ5H9LqZGr6fS7
EabeQglpsNsS2FCYBvtASSGUl/wCBzuvavz7zn40SWpOKmqN6Vk+mZXLJn+u36O2
Q4FL7CAv756qdj0mDjYLE3XmE4Rr0c10htVPEQlcoxg=
`pragma protect end_protected
