// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:06 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UnRHvSk+q++VIozEFYCRu4uuUZD9gafPA27yS1d/HEMg1vIFzj/RfZGzJAC3S0F5
VOhbPt4IssV/+Ux0oB+YWp+9Dpl81Pgpcmj9bqbKB9Uq9ABMMIBHWeOOdoORqLio
Tum8GfL5K8OTZl+acnrnmMiSqoodTyrHuYocLSw1fBA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20992)
/ADWTajKaXfQOb672LVfw+/G+eIkkb24Kqt7Go6nneQnmbyLmiPGmxB3YvR+OWLV
q8z7DFtebytZBhDG5sN1cVa+76AgopXROq5txbEBcvbnJnhJihGAUng/UGZEbnKA
tqtpnW77NtZvkm+DuPCd9NTKqJGDPgGag/uosc9cF78/Ou1Q20sn6mCiKFk39FaE
TjeuDvKx0BGHKQiNQ6Cncjr1rab49G0yoYRNJV/Ziw+uNKMEn4vVHE5aAU65QgRV
T+4WeEwLnTaS38WaU9vluwto/JvTyGFgz8UfqKtDQ7rc/HtMCnhZXt/i7bID03VM
xoS4hAYBlWVUvRy/oo9l+dRIKkCoPvrCoQWfmTiAfAmMejhqnJH2z0HGVlEEE+zT
i1HHcjrFnmEo/Ti2jkMKDT2b45t1KvPdT6TQWY7LWg2FCWlMamguxhbS5rSHPB5F
uo2YtjEcxIp99UCqHHPsOYXUf/Cci6OiHXFaEd0+IP2fXq4I6Mflaw7kycosFjCq
FLke4BXXbQbhds5x9ybjNjEbTcnvm1Hh1e2WqiVaulhMya4kV5Hb4qRhiBtYTn/2
sU7CL2BtnRz6tAF/rp4liDpdsLQ/W6isQ9nezoYjp1yGwSY0APM700qWL/eZWpfR
foVmTdc1lnIhBW5qDqLUceU5ANpltDWKZfrtPI7PMX8KPmjzu+z2ofKuF5v/ZXV7
+hYy0nwnhKKu6DuxxPnCA8gkVqV2cj+bVfrBHGI2Xo8+B12n4L7AqkaWxlwDasu4
BJI20YvWmVWPs6i1cqqi4JCGT9HhEwiEYTUgt7jI4YeWbpL6GpXt+GfPQfDop9pZ
v6OYBA+jYVjJBMyPMGueDEnXU4LHidd9kE7LbqmgDKZfwo8G+DZxjD7enIlQzd4P
GE9v45hNtTFLacdZrChhHE4C6zD6wlqkgrBF5jfP4DePrlOl1Ywj4cfhSm50Yvks
eTQKnTeqLJ2ajrXadzlFkQ9hHyWko3xRMIRX7qq3iLuWhohlOe301zgo6Hs7F2Cd
3J3TQIUcW/tHXRUDlMT4Q0ZY8Rw0e2gUKFIQXbnTuX9WFRRcwwj3wb4N3D/lVp1M
YfKG0ojd4iFLC/gRZhnzHv3GxLPGQpQhdAukirBkJsV2x1Lg86HQKqIc8HtL5N3x
t5nPn8CAmihJ4Kg+QCGUPipJ4gA+MKF/+HblAbw2aKAx/OqhJB9hrb4OGUIPq7CN
Ux648NhwYxe23gk768RAEAVvcTHmtHQa4s0b8dyu+TIwdC56q4hxgfMkcISrG1hb
Ht2HrC2Z+tuvXIi+t6+/9D9HIdvdyCDU4vzAPdlkrSagiMAKGarrQmm9WiJjDfL/
bTiFrA0ZV0hYl/kJTvhs3fY3iugLmXdzzjqZLU9LteHfhChm1UxSIFdzLQh0wAWO
fsXEWOD8VLjfy1AUeqQqDqzHtF2jCStqpwqIMgFm4oRchGpWwc8Ef8LMDjMi/KrS
mfKLYwO5OwxqTtvoMlbkEieeaBSnZRXRKWWCOK/FXh9CeszmZ8agXHaIOv9vOxFK
/wiEnt6zujdWjQ7rslkY0lhezZH+h2qcUwOO6rsJuzOeM084nXz68AvJCP3M5q+2
gmjJgCXZV4PnyndVOF+kSzsMMuIwbs4tOyaOvL4DAbnwM62cEd3jCD2S+2KLWVt4
vLnFl8xEAC1ovLoW97s1i43E5D7vd30OhpjONcYp5FDDVv4f2mFkII80qGmls8Oa
wCmZZuHgOaYP+JajsACYHokceJjTZy8zZpOy8wpE+wy6/L7Yc+VBWk8xAfZ5Mi0F
QS447GHA+i+BKmuImwLiJncZ0KrOXSMO3LJ47KBuf1wuy0yUgbB02O7wrFBlmS4B
2shg7pEcBIcYarBbWNcpAWlsXSDouTLoUsPi1U71hjoSr2eemQMZ9SkAqObhMM1t
AE80tXMzUPWImMmq5rpBQ+s5y/5O6jTF6pWrulyua7lJ6LP4+pZ5kf33LwPFp2DN
19UkDRm8BXfOABABKzc6vASynVTr5d937DcojKl2p2tYemHet4hStWs626l9VThF
eU36GzorucJqxvEuMDx5Pa/UjdSeyFGyyOgPxxhyc1eSoBCKm0nsz7zyJWDUk46a
GlSJ9Bv0qF5Br1KwLZQsmhzEjPlRCIZoaLBoJN+PCcUiQAd0PR9OYvlrWSncI1wW
3Fc0/b4i+GkxB8z47eN8E/DbIx/mvvStpIugGXouKq4Cq0JF/RYd+ySA2sy4YISF
Rmx6p6Hw3uE2F5MzyYL9VPF/y7gDF4elF6gfF9hHlwPhcCO4UviY0sH0S9PmNTs1
u1Nzs1ql9IA9CrOT76UjrJ0jkrWl03jFNoSL3fCepY/gvGhHCf9lgtsuhzQhvLpP
y/JdLSm+orbIrYjxhcDX6HC2z7m6eeA1y7p3DO/hJxbfgnHRsLwCu9K6EetiDGtY
1fBnBf3SmtBlbqUlRbxlJZmGWgs7NKEYTrvuBnbTvG0NdOaDcY7wtFvRrqcWPnSN
ZYLWlLQenf35RLw5oIYOfbTyYETp8On1xk8rcTmmHDa1MZiuVSBL7wn1T2u/UODB
0hQvNlBdhV3EBIJg8D3Ft8IDVqxBpl/+PZD606vnx6e6WliOg/St+NaQYE0K7gDm
X70k13mYofgQNGKG4jpluRsv2gy1RlcNmFf5rXSYrLtk4xAMRgzBYqbPVp+k5cdI
v0v7UipaQ3Nhw+Qw034SLlmE144rtX2gkAulCsvetdbLnJX4AT4T3Ce148xOE1Lp
kQQKS5QoqcyWQDYcFhTyGUnch4vsmAzjPLdINxWlLlWQ7HD7nm36I9EG8oShbw1U
qJyx1BPoqE4LC1bBP7YMPgLFRcpGYQY2IjqB+ji6QbWzDDoumOxQfduqYjfE+ffc
gmf+gHX/ev5Sulb6uOA9MzaDkEh5ftIdcJh2ZcIhwOYi1dVVwmq4An2Eih3tG2Ab
IrTr/YL7BA6YL8xRZlaEJ+YKxXp7Uwy417vabcG2tlTD1bPFpgTmjTqFSbXugWs8
nHQFmCvM5/IJx01+tQyGo6WK60BF0zgCvq745Dxx7Z0JR/C8DVLfmWxsl8SFcUQP
DLiEkUnvE3X4BxxrHXO3HmAjhBbhI+Qni6SydfQVzbjysAAjb8WBHG+nl0GyIpa2
F2NmEnMCl+LBdBkAVtTiS3aFG1MzEHYJjvdAwvzC8elPXCqZmbjfmfhybUDiIyM5
yWJQd4dHw+O08qWoUnsBb50GEYAukInN9DDvJeHUViibluL7dYT+LiVTjN0SjCMb
jRt5y0aevUMvrKsXZ2jULNfMV0UyeR3CQMjuajE6kwHAufKFZJPRKo8zv3DL8brs
7ayQnMaXNrVfyDY97vnb4q+RQaTCZI7b/UYfBKkGsVCwGRy0DcOp+dUtMnOfBbDI
Mu+Kvqz84xhWwQIJ7/l1bvQbwu8hHCyqik0rm6jGQ/p/KT+rEANb/Sen5YZQzr/x
jRxFWEPmObfFJYmt6FZYt9bsd3tFs+SwzbKw0MJLkorJNKwhW1jEDGegnHsYxUQW
z2kYOlNdciCjhu7oKZPPCXZ+GLnoOw2z/oUmeBG4lVaJ54iL+vK/m/QO6C5S19WI
ngB2+ji+b9ZjM5YOqiRSA8gykp37MBi37BY5RJVp2pFLSF90m5WaritS9/t+CqGB
4gTzGBbxLFThlLPeYZKALeEd1Fztk2cY+apZAyFmiRKKeJdn/tiH9yV18fYO4TXZ
Um9v1ptv8MTCKZfJyCDhwDhwgL52pcMfHBzKrxmJqwSLp00un+WA3Cy14lrcfMhE
L3V7+wE5fvAzSDAJPnC1KKmRgXMoVoOW36vQtxap+DxMqUEi1DkNJd87wmKl7rkD
gqJSFfqcO9t95vnmkPTOstM4ZD4x9F+61H4VKuxZkf/NLkMI6V2GxHwYjCq0oGlQ
N32tI/gWYtbn9qgnpQzpZFxsaRk/FkrB5v0aOFQq5OQTtxNgqL8ceOc01R7eKiCc
XCBechTBbCaihrjKEuQ0QqGyMsoWOLy26Anz0XaozPdruZBjw3q8QCatKhdKgaZl
W3EVweTvC11UFdtBzxPWV44ouLVMJf0zZUgdenuQzZVkkI0Bs36ITvTNdfIPMIw+
BeuMtL+sM9AWQ8ZRhsIxGHgUqba6ShNpbT6JjTs9I2Z7sEn/FArUcgvj65m+ZK9H
IWrtOHyYX00SbLNiLXkUBGb8/YDTRAnSHC7F9xAS1l/8EQF8CkMltc9AoTX9Uxfc
lcTpgurqcVQBcfTNB4Is1HfoviBYvTgtdyNQCEjWwvhDbT1MlIQVEr6RhEmZtZiF
xA3Unvc9ruMNOxR/FKn7GyXAoSJmKfdM7ZY+9v3m4ULBuPNMT2dInVzqDNK3XXzX
T3riBxzDvsrxQBIMM4Z20s2WKCIZtyyu9RKNMFJQC9ZJMVMX17mHsOCcF5SND4tL
4LtFGpmBL14hPEK466ay/JqtUh6QKTLpsTn6YaVS7kag6ty+BB5HPmmewQb5rVfi
nOwRqabbtvMu4IKOwkQ2vMvoXjEzV8DG0J27U26qRkH7gGRqdJElD7KwX/gq9MhM
iWZqiSEPxuTTDTrOVmipZNBBE8tzy977rDX7CBvGXYUJS6RcNtKvJw8WwNnryvMV
uiWH1L56hlNuFJmlDNoipZr6RxWEN6AZZjVr2pGdOJcaXvf7JGTDArpXLK/WiKrM
+E8GZwgpJKkhO3RbziETvKfZoPUM4v4f5WNryjDe5cM+ZaumR9COhIIQhlMN6t83
ZjGpdtg/6zolPzc3IgCGxOSpnR9+oiZD0TO5PkZnI1j5QHQyyGbFvPFKhYgJMS7H
O8Ake5WkuVUgjZHfJ85cquVzgzTmryZi5faw7P5e1ieV7HbXOtIul9TLW8FeNDck
Bou8LrLnwYpsVdL528fKztFbWuJULhQ2x6Y/yOf0sl/bigYmePtS4fTQcix26GTS
iSfklLr45lMno1Kh73/mMp9mog6HT3gCWRtwZ5Q/XlQ3VakxEn0mN0GaVwXZUcn6
BF4uvdlvfQ4DTrRHWq1cB5GWaw2Hs7y3w9MsQpJfnoN5bCGjHG05W8h2nzXxsh8R
RSk7HlX/LKE/Jmm3O1xnGacJcLEGRqGbraesnOAyL7z+lOeZw6bSFaghl9uZMIVJ
E78pva5OUgcGhrQIMi4d6y+cBrvkUhbo0j2JbjZ5CM9pfBrw64Y9RzqJSUjuS0eo
wiRjR9jZzRBviHgNmI82JDbnTCkf+O8Cxdapzs2A21L9tv0Kx7TC+T72H3TPOIv/
sQu7ilvERymQHv8kgZHZ3N+F9L0n19jWkhz5p3mI8GOj/GZsHjl3moMaEv93rssh
mrTCuytstCaBgthW2sHdRXyNSUCi4ZfxzUWKeBpFhQgtBnC3oDceaAYe5mqntlHc
vVSeGYmZkmi3Ix7nw0PxCgWpBZ/ZVRklSCYmWHdD7s7SBJeVukM3jrngFCcTPazG
mkiL02k3BLLbu+i7T2C4zGyLbEt+qb/ufyjz+5SxYq13Z245QZs5xbM5OV8NS7iv
KOKHrAE0apDmgN5cf+Pf5bRiAc2ck+6vwgfELYTv3K4IJ2Uo+tEV7o/vhbrNcjLH
6THxHSA+ayl+fVgNiZXQqmWbWd2q68mzz7ziheTQB76svwLh13uQlbI1vDNnhpga
VE1WJKkbkXrka5C53X6QUVorl2DyeEmSZorRfT5FXP1Qy15I2JstFMj9lWnzIQUN
2JfgL3Wq7fnKpBvq16b9V3WPcfNhW6GN5aZwAypKRN0pxnosN7gP5YCc3ZpKNQJ+
xzzqtn4gbXUbnFRpD4esAJ4yt2j8fuVKQdmfRH5a/wcuwxqVYw+SAcRSYUYjbK8t
Uyn+uKnabglk3Gpu2DB4SHCjLOtpnEOVqS6LXoetuKq/meyqLgXs8bDOxOTKXSJm
uUmhikkLpp9WZr9QM+e7XodIgcCFs/y6QruaoklfVYrTyfxqbesLBer/MtbMNno9
8ZNKgmIGuqQaTxn/nnR9DrohPnWkvlgGE5hGrywa7qpHgaZxZtzZezh2MCHYM0Jv
+i5CnNiVI9w/CN6GbhjKXzRepm8wHKkxk1xRhtEfXZ/aN5HqGR2RlLAzWppcr9Q6
vunBYm16emam3xygR1eTKFWNGsf7RnHZEawFEeNwGsMsiYmVBElT7/HfarrfAokr
KAhagH1kQsGHOIrzy9lOvtLACIXKR6s1/mgwVWE6W+eCnLlKKE4tsQTOn9fx3gYE
rto2crgWycYeDlg/l1sg+LcyOD12KsBc/CLpnxnH8UMj3kua5+q08pi1eelh9OQN
a3j/jspdSyzfx0FhSc9s/Gi7tmFkZLBEsknTR0Q75mrmyZPpYAcl1Mxk+mfYUQdr
tBMMx3Zqt0cpRw81aBn96E7oI0bZxYhH+sjO6zi1iew/pI/LOZaxjiHe/0dnUaNY
4B2zXwcHksI+rAxCcmgCA7C8n6oNvlnbt3owwJUtr1+MGUMLiKoxbR6Fvd2d/0tB
Or127bamE2HOpCFvZjCYSI7F08xYtmAkqpGWef7ccn4240f3lAzC85iw049Sraiz
ZaZ6/VBLgEqYhJtOrcMC0Cz1gn9GazVWI3BrYSho22Abblr8ZqbIQNgqvNlVhykg
mWjTUkwBeViydfWo9xcAPDVCltriT+ovqTHlZtSv69C4FZPj+N14+4eeB4mWrJBd
fg3tYm9DsGlKIjfJjusA0jGOXcPjxguAWAfB/se63F5LVpmzqlTEp2t6sqnSHqRs
HG7dyQtPxkrQzN8IwRHhYtO1xxVWXJvhNStCMFZFY93zWaMSDCTCoYtZIj1+Yv/k
jEF4U7OvsfyP1ZtZhVGglIKvpD0gyFwoNiQzZck9pi0dZsHCsEGtQ4+VMePdh7r1
zRXAHAFnSCsuq3K8XykmVUk9Ag3IIkAfhMtW+mfIs5/0UEOmUV911tmpfLE/iSkF
K3xLcMHcjxOwoh+inTcLbsFWry8oDb7ODUqSA7Qc/tbhdc9Gc28zaAzrBkF4XCgY
SOvoW9trqV1WVAOAp2ALXIuChqe0tyL/ejZdi0L8Qc6rWnrH6JQWd3j2Miv85RKm
Cu1+JHKFnaBKA17C/Cq/HDU+xlyg3/SlEd2fb2Y/bTMxjwRMiiDGTxrKmG2eflz7
/nmSd7PO/lUbOj5eoUVuMTMF11nOP60dWHDHmZ6+Ydp5kmgIqF93oCRUE1wMpAcx
QyljR5ZEFB2ypeWWftmEdvQmgbqXWpVlNMvVi36G/+UhmlFxl0np76g8DP+O5i3Q
9aFCssAsvlmSvAVeuTGHYJKuGHkhMfe3XlZXmGMv7uk+1jCckwZ++V6I/h2PU3I7
gITNYTrU3QVXg40jZ867lLNK1PksHeYrJB59ipXvA4+hFHxWAnf+Yb/EsUX3x4iY
QKgiPy/elIEr6FarsNm9dec1CILI9XZzXiWaPgwWyNNbKEkX6kxNyncn0MkqTcg3
mM0ej8AJWEjqRclCwbZbRPM0Tf5kZSB8t/SlQPMOU88rkW7yuGsAQbFFRUsqXb/g
IioPN4YpmSX53C18NmrQV/xsvOdLS0vrkBIcExbFvcI03uJwXDnTXlA+ku1LLCA2
P9zS4RLFhfaL11FN1fdcDy4ul1K8ocYGkck0V4Drcq0OlWSMJsqJ6BYzQe8RGMZt
zh7Hhn3EkS7vsPyTnRFs0VvI9hLnZQYU68yqhYuqYD6JhXPJk7N4O3dCWi84DifF
c6ns0KTiKl5/jikRWhW2qqGUlJMdObuPPkPgxcssEydY58NvnDL0m0/p9vIWXRFu
es1P6pYHa8gJnbITuQX/PaV6vxwhyPhqQcM4K9RaHysDz9muRkwCoBVmupGy/GUf
/W2mPOXBrxpVVdxFxQ/mYX5fIi/8VFsYMOfwFUPwmRCqLHsxsPX3uVtWirQqY8nq
typy5FTS3a2O7fVGsf/Y7v5NA4ioVi1GDp7MX7Nu3EG9HTZLM2Ra39prdny5+MGw
SLv7AuO+mJzrYxP0Mkhsp6KdfqYb7WNyMqbUdTasnXr/NTGqXctbuAMFw672oOdl
Zyo6BQnqp6rwMxm/QRIVMX9d64Yh+aEarDHD6HG8A/VnHLeG7cU8BdKEkYIZbLue
2RjK4lBV3wyfhpgVOWGdNaMe66AYSK7ugKAlwH1ARmlTBHvXSVts9fEMMZPyBUoy
PQuJwWVwVzhbIIKFigEo+Lg8fXQ8AH/CV5C+i/S6sKIuoStFnCw0JA+kNojNanvw
g7Qud+p4J1FIzw9qW63D/xekh22QbiJnyIFqPd3K43+NrfBmdJEPSWrRqoyTsUS0
AidbpEVzRBJvCAyx4XfBNMn28BfrbZpW8SiwJQfrKZF6Y/Hx3DnJdrtrIzzqHkj6
fic7U/XjoTwySMtv5iu/4h1/akfeU8MygEPCnrz90vPcJwNpKkB6YL6aO6DIT48h
64OQ1vkQXRc9cpCd7z8k2NJ1UPGot6duEtEtJTx6dhkiwtc/azeCguZl18yBoSaL
Yajrpz7ZFIK23S3NIVizfyS1NhoAhq4ZCijT5cB2HK1E5lgLJiUB5CVuafE8DeUz
j6I4EThwDNxgTBFsgQzYnBtiSnopdoGhpd9wyL57dajYdGdXXLKwroGw06jVk2gP
MnZd6UIK2BusVuc0OcI2bzSe1MJA0+J2eYgprF0GkPEOp+NTEn2RVVxaugcGlyvr
OpzDrqUVowwMFDVKS8gY3928FRSe86WMyS1YPosl63KiufR9SKaZrZk5dRyvegMC
7EjyPcY+Dq/0rzRcJH6lPQ6SlMisv8FWOpO+Ftr/AREapcCcdlmIe3yL3o0ifQV0
fg8V5CIEDDdRoikEoxRzcYI97kjFIYVHZgu3KHUX4xlmyDDOMR8820/XZ2o44a6d
tpVdNwTq4Z1o+Hn/M4JZb+i24QE51DNm3yBVhbfMNqV4Hd5DBuU2wRhBBGybasDR
L2DVQ6J/W6/KKxrZ7ahZGpqps5Mt9KLR1Uv5J/qlbTERgMXmDEgaG8ymiIgaIu0q
YsNqV4Tejd6hN/A/lMKAJjztOBEUQwiHG+ifJv/lneQnRX/VbeOdvUHZs5TN733H
Yq/DIsW/LtqwpWraHdUQodD7k2ANaVIK3bHCoaZA98Q+AhKeHzTtqEdC/WaTnP0Z
Cu72QYpKERNcXNHfnxEIJ9r4BFNyAx3h32dtKOB8GIs89ovXiZ8dRgzloM5noLBK
nqeydKRR2V1w9/BuYMPclmM6RKDGcqEepdYFXOvDUFndD5Hva60XBW8M5CZ7NcSJ
991PiUuWGLzad3cgrEhMrSAw2B1MQmYRea65wmQLrcGkO0gymhMzsVSXnRcAHW3J
2k6eMN8Fa1ZiDSwOP1ToOY/8+/ZdyJzjZ2YE0MvuvVcyFZR37wts4cqVvIzZikKZ
0Q/ozy3mHV/BUkfLrALwMXdFn+GD6KjOwirIYuJsNxL7G7pmu8UNrdJtThnnsZqk
VgdjdAM+xouXk6Nny5iZybQOcN5pkV8YtCjJv78xnIqFepqHldm6eTKBndHkG3Ck
ZdMnmIJ6ulyb/Fst9Z5/3WGgbIH1+9tukU0X0jNuZwmlauEiB6Mnv11fxI4uTnX0
b/gLsitMo0GUjK/GSJ2EvTsO2b2Kx7JU3cJA9TC9WCOglNP9hX3U41OwxDy7ypp9
5ZQAkuWyZnrml+wgGedjtOH/DxKlFjy8GNFCl6zw+NLDzivNWbrU2Rzj8LSDnhsH
2sXGV2hsW51pQkuA03sOrVwbfcZZoDGl/xMTCkoYRMQfhTs8AT6DnqjqbGhALj8a
u8B2S9dYQZ+2ve7pPl+AdqzT9w/JIH8IbdyApPgxXCTUnwZzIJY2uIjs3oOQ4VFA
fyFvUCxdhkBsy6ZljbNRAKYn57YFQCjyDYKDVK4D38K/xlMtH4SqVXpN/lrXxbhb
4LKmqS5pNY1Wvqg5jzE/tZ3igSjKdZTBDWVH7BJo3vKpbYsRkmF+RZKnyyDGaqHv
LG3E46A1apLkQkjyg05rLnJzITQsf8G5vNuWeIWSnpNuIlXFp01OIqHrjcmRtr1A
l0PZyzdh5hIhMK2PsZ4ptP3+WRI8VgRIQ5U14zLqGVzseAUI+Q6om3tlW0wJagpy
Typkve7it3zdJ7WBMtCTTiSl+QDof3pVIVoEkM7snnsrB5zBUNGkKy9Z5OaIi7eb
mtZjKM10X76zxCErwdA+DoTDNRW1jxLN7pwRNUVZZzf4EwJwZb+1T2IBpURaBEk4
UB3Nopbf8DDO9x5JQMM3ZZmFTLH5B+24jvJIUBqMdEWBLtbYFWTiaydUoukakydG
KgiiTA7q3KHQwKkNgx9rwutbLmhpYHOuBEcwEQpCSqGA04TvCD4/ClcCDIZO9qg+
pl3APK5fAkt8T4v+vuypi7braOI50MdencrL1GplCk4K/1KOOlWIGT2pLmjErtem
0pq9XW8pXmGMh1rrWcDiipFuc5qC7P8JalkgbPQmSfHeudAJAIOQfNO35aKKDAzg
2kFUUM9zsE6vem4eI9WUU904qswCNpNRKC0qjmEOfKWcjC8dlfIc2SaZie9d6KlL
xhvgvYI0bdqSG6sUha1d+CpEOY6u42NAFVwkGNOEENPRi9Lkjw4UUs/JuPJ2lOPL
SFaMWsD/dG1nGExXF1ylYiNNBjGg6wgeHHcTmlkUbrkPFRgS/6+BD16O/oJiTokf
zGeVo5VD5RX2LhoJYMr5klquv37sw91L8kixXewlf+zNdR2VaMyqKx090XzAt7zK
e/wUtZ0WMqGvFMParq+mV/ziiJZsk8eWhGhXFtTLT/jWEId+9RijohN+KN+aQSpw
fUKKLIR+NlVACBLbpxdP0oj41a32uZHtYtMr+EOhLJL3aH3Moz5ybFQKg/M9w9pn
o5z/+VrHifNV5b2uGHXbvhfAcxCarBiRX/rHn4v9UMKw70JoHW4vp7vYdd5cbWrb
1MDSeD4d72suraJxFAjnFuDyhbhOqZee5DhHrmJM9M1Uo2HWqI9p8uDZ3REfYfjR
epu8Cs/lnV80DU+5qj+lhR98Pp4BzcRCdBt7ha0krhjzEkqcuspGgeFUcUf/eapK
YAAvhHcCJdEzi/9llXe52Mke0mU+E6bK79qBXL7S56DNgaLepq8gZ9j1S4rs/+H+
ZT3L3Q7jfdfKoWpag7Lw5Sys+X9/TtrP9fbz1MIV5SD8k4zFjMmou2/vfXHWzb+D
p9iRpP5SKrUBhfq1zV3V+jlD1MbrvY2JmXZ4JU9Aq9jkCv7/eYWpwPH3QVvvYOh7
NHUSilFJp32gajsh+fwWu58OS+yyS7bfjsOPCm378dCm6P7OSeSwzplwFJoMf23t
jZZpSTf/NyuAIXKaQpul5qIYOryAs7zByOPISnEW58cVPBOx35XGz4eN72fYonle
Ky+XXsEN2Suo7+tt2YjLdYw0R8kL2Soq0YZNv4zQyQEGt6hAYLP6LkvHHmP1uIir
rO+110MMfgeTiu8NDdt8xG90SAmt5lMHX5ljLxnkHOXJyi2TM5IlNn/el1EHpboE
Ebvuv0jPKX7YmiQAzw4RunN/GyH33BC9bGwmQYts9axCXWxHsaKRbLUz5U3OB2Uc
4Md11pIWWPveP+ln3gyUQT/aAjpAyoWZYGVDkC69l4WlesQ8X4G/2/Vk6Ehs1KhN
xSVoCTkjqhABTmWYmUqH05NSuSqQoLEC9eKJUQLoroO6RVEoVbiP9jbl2BLvl6vQ
xVweB24ImPVEw1+WwIg2VaKuMx8XSK/ZhKXy/caaWwqrE0TtNJwHyV6JRcPLT2gX
UyQuRfrEsq9mJO5zM0dDhoneiNQK9PLQd5ZM+BUDqZxEMnmZo5CxQfnoaMBhynqu
eSv/JThsVG6OrKPdtVXT5sy2BvX/ljGTMVnyw8Ntum4m0tHE1n4FvGyTCT7Av+NA
IhQ61HW2xioWcplecQDzZinBGTSGZLn47B5HGXW61Xpmb8BYjVjHY5fopI/1fAfE
6PLgjRzTcqEpLb6vBn5Ysv1THS/oktmcvjUpEl5sX5O+UHP/NTGQJA2Q4BQX8bYD
UtQOSjVxjDe8p/ML/n7KPlRAlUvP2RZzf60fkX0is8xb3SvqsJhxGeejZJQDS33K
UjVxbA8olOkaSnRyedFVkmbdB09fr0uFDnIWVH5v6KoivAmyb/jK4aVTY2l1CmQ/
km9uEaBONw/BfKd7E0bSwR3m1HmgsEZkmbV1YOrRgsJIWfcc/jM0U9jCx9HrB759
Ql1QaD1aBsZpuFNBQhjbmshoap4KtRARHQJYW977Am+2gGEjZ2L4SxJTTK1BHJ/S
4oLjRED7fY0zIERA2oV+FKtLBduSpJT7EWix45hiSZpfFBZxOWZVDfO0Yis+4o6c
FwucypwJQSJ07fs0iHlis/MYcWxQFXkpzA2/ueJxMjO6xHhAyx5tYpTyD/V01lbD
jRIXx7/DMn/NRvhaJAXudCWMYmwiBbUW/tecazYj2AZzYInLi+/wAqQfqxfHs1VN
6VL8hiT0JuybsXGBVCVWJiKi7ZpqTPxR1NDpcYFIc1Y2vBhv/KJqfrl2iKLVnike
2uczU/v0AGlGc6pBKYsy7WpXUgwGqKwwEn/FMFNOEE/CVlAVfMmVmlu/hstJkY/k
2A9EYr16ens1SQHqaMGmgpy9dMnH6T/jGFQ43uX+QJiHDWL1jzEtU+sPvXyuoXCR
0feE4RQaPQVKI3/LIoma0GCUfD6NzgZ2kFm3wydLoCGrZxtWM+8g0xc8o+DpOuxQ
5sBLeWY2HMyKGM1GubUlLj/w6JSvPFoNuvWHU/2KUzTmVjumYJVcHaDxrglMtGmI
QQzBNgxopupigoKqYgJiOrGPVgAsqTk9aviVoPBl7+8GDylodMZWLhznHWIgiX3f
KXl6mdLNZ36OQp6Dtorli9kvBEeSZyTerwPb0qBGuwPOjJdV8UmeJlVd3HBwRemD
gVK9rchNMsJFLJYMVyjTMyxaz2GHF+I3b/e6SX9ZjK0V2KH+dCu6XkBs7dGgfObe
gLBM5QsHOxdObOdLpjnM7w7O5iCgloIIKfzlDIkBZhwR4jurJBx2g2poWixcpOuD
bKWn5fAMPBIfUodcJMDywidkg+AJ+4ASrc0BgrEY7x93rdPiNCc75kr+prmnwU0D
8ciXvo8h0hFyDk7l8JHgQ3+pYC9f/oCZ4bGsp/pzHfbP5BqfaNTMjOfn2EpEtvtL
68Iohz4sPtUUHCMfsTmKCAQ62jYZW30eVORl3e4ne/Ipw8cSExTrLU4yKUbnG0r1
haRP3WlXj7EAf3bq140kPVrTfLM+GT/raFKKupbLFBr0dU7HKVEI708GotgofTdi
bRsaMGduAFUw1zjd2ldA+1ujViFDAnqbAfLuwR/okta7dp8ZmbMKrp74nLL/596S
qrQQaJA+7fsAsNvJ+X4zb+HkpMxteCOXimo0j9lQW2Wm97ImtE5tipg1RzhcdG3o
qnm8bPekKYS/goyjvF4cnv6DTfUI2nY8tMBJ0uCLGl/B8L39CC7LEq/vNL7tnHMa
kwR4RnnWUnvrBjoDlG5b0HGqRSJuOddlu6RvbVWe7LhoK2nKGck+PT4yg9rNFWNu
kbqn/NXD4oTnXbIg1ye9+V1hnR9TP35sfq7EBEzo3VIE8+KwERoLBlsQLW3NP9FA
kJ6fyvrybHrH2j6lhlJiXriDWj6Q6Z7COA1aQDDkkYyuLMmVCKRBnVaBtoXaz5fS
+lQqGGJ8aYpVYcJgYiNjwItP7YuEKw0cKeNFrM94r+6KxqJfQza8vxDUug4oI7Uu
uzIJU8+536eG6CwwXLhi5sCxnGWvmD5QxW3maFBFNBdrqpQrfd3hUqv81dt6Zcqb
vF9NmHxHDTlpVNZTnMKzVlzS5hn/2SolsEFTYzDJG60SmYBcf+hPByPKR8pWixlk
1galVcOWWMshm1EvzHwy1r+yVSa2SR2eCtFCDq5dyz+Z7eS6o+CaLFMrQ5znVR7u
ar+fcblnv9FG4nHtwGRO0Qaue0anA9e1i8ZKaZRxTxHHv5GUcXCPvHndQn4DUVs1
OrQbs5v5g8nHmd/ri6GUEYFN94t25shZKYBftGKPxTW2XpgozSLG5uoGtSpEW67M
5Hdp02wGFO8fYy+QsioKTrkwRMQDGPGbmq0WKpriiHwgRyC1vRSz0dQJVgoBlzTa
1Xk7JB8YRGOrj9DSM4T3P2TTbZmQjjRFND208M5xa4+P7Yc34d1NXXmVloSdW2jn
W4nisyqOZeuUTHr46ffa+45/ghLWIbyFIAt8gaIr9ksEnuQQ1F/gqZpD/1I9ZFOv
93nMpqxrRwaQ9Di6HSGsgrua1zajX5gHQv9t6xnWugjFf9GXrOl0SKDmD8c4voBb
hQNSm0HNVvANjxeDB7YwGRGg6jE4vzyByLFx9oNDdbdqoVC6gLZlq6iYdRU6tuZv
s+2ch/2H40Mwyxk7zmh270q2PYI5nXervTx0uE793DP1/SkwaJDks8kcltntZZJx
mEccgn0+7onnT6fYVMZ3Y5CYS9D/1RSZQoAD+Z2fbHRqmJHWH0WminGdUO1w7T+R
25uCsYazU0b/0T435I5X3NpEjyNzmdZS7m8r2Lf8MsWJ2UQev6ANjZj7I4QUj6Jh
90U+ujUEiwqj6NnNor0qfsPJqHFVPNOoQyXfOl3KbaRUKWIrrto8LBe0HpJjWlNV
x6uBrShz/TMMW5Rd2nhy4QbX8AMgUe+zwOzz71LMrceoBjFygKDId6lqRaWltrnC
K0Sk2mNKE6tLFRM0RUhbWUN3C3/t6ssWEQxJkofgNY8P9Pg/hftjLVk/OtNmtQQW
1bzahcLOgngkiEGFsRV3K9CYJchX4QnAbw45XCTSvBMXY6vVb8jC87lrNoq8eq0/
x5DXHvBrHfNG6drCzMbmeP+fUkfx9RinhNTzlNWAyhIhYH53XH28IJOL6BeM0yjt
uCBtjRptsK/zh1FXZjbiaJQ7IU0xjwTCLhXlZ+6mkVddSUydfsS3HOY6cpWWA1B8
EvYj3AV3spMq4PHL7AGw3MDKQOY6NvLxN6ynefdO1aEW3XiamNko+JwKAqmP49T7
hMADq1MPYdf36BeWBq/gS/wpFGa0q7gZ2L9g9HqyHnjjdG1JcsM873NLnxyOGFgh
6KoiU2V4E2ZR/8F8L7ZRfF42iyclBVcLkOQyxPG7VMAP9LbRc7OzSd8p9kXGDI1n
N8+PHlXWFQi0vZo8WljgBaUUnOikwT3g09Pa8H6vNlBd+zqfRH2st6nfcRqAiFWc
1f9O+mSvtWkTmh/3+n8rTAiL0P52lFp9iszRx5eqpwyFjZHBc2ItwBynNzmz4l6X
F69XHHU07NYzS20zQuoaHwsDvKi+nL0W6XQbgAM4zkLQuGxQoFNN1n7g4/kE0363
+ql2TCo/pfmoilp8hQSluRUI+YrMXos0XHIF2Y96Q+7N1VKMavxrcGsapavLue9V
xuEtzJY9JMtmiwaL7/4DpBvQUcO8ok1k1tgGI74wNk96TP7bpjUQb+p41BRtza18
6rbvjid54OsMZYI/n5bZ4GCVj0Qd+UNN7t0z/6PCZXv3TTVfF3ucSa+jHa96gK+L
GAKVdeZ5m60GkWP6+ClWZH/aQ4DpNU/gnm+x/E8cRd5iWXk9L3oEM7lgXurre7+P
nGY15V9ET4+ExMAeI6Wdid+SFf/0pbaALz9gCUC3ThS4pwLUSIf75nK7nLOFPXe9
TnHXc3B4gUeZNTH/8tddW2jAi1bfaCeAS7kBMBqZ0Uy190LpCGhEl0rXAMXxEVtT
TBarz2/7+iEwrc4Z5nue8DvDVtwZYXsTFvkzjb5Ob5C2aCExVZ69SWgpoiDJdndc
+w80hTObkQSgyuaAgKqWKM5lanp1sAKpI+M4yIOoSbd3UltvoocURIAqeeXuGpvS
kgYnZC1UWKgGXIRujRQwkqpXQjIDvIwVcWo+bO8NDrtKwH0mihibSnGElsm4smjb
pfkANKj1AGtUet0aAEg9fyjohcbOr4F9i661dvEbJNzy4gZxHG53wp9pI8Qb4g0W
yTrZxJ0uUbm3r0eFCknSo3RaTGzcZ57wTEMspZPM92ZdvgrjpNvhxj7D0kY4Ji44
rdN5u2deO/hi4yKwU0MHXuc1iWjbrAXwghHtkEn7GfVp0V8Ur/AJqZikEmQTRQp5
wvHLjC2dT/6vQXjNH1gjDo+TskDxJ+SlXnUn5B3wlc2uTcvEUD/Jxpf9rhSlTlvY
1mpQkv0AGK8ghFjmVk4fvzeZECTBSYjfcCRdlta4FyY67340lyxRhbVGcARDl0fR
k5qv0GmsvmoHjBG7UXg6NF5kqNaFJPqG8rvUMv4ZcNSvOLIM3mUUKaEKKZV9vV61
ZGcj8A7mE7Jd5NYdXniV9PbdooAD303HSOMSUxSqTE5uKa10k30dW77PQ9SnhhgX
dl5QUferUUoi3eqHdMvs4wvLLQf0J60/A2LnbG1SoVXQlPoIRJ/+pUoZqbg48Ggp
lzDq/e4UsP/Zq9f3VOVeSxEZeoBLHO1I5OABjt2SEauCIQOUvfrdq7UQurto/ZL1
FOlBvkc0hmDXnnUPUyUOi0e5e+dllZQhTB8le6viHF4XcZPt24Yo0AJSB6qD9A3P
M62zG5BrHA5XGfbH+/OaNehwTeqAoJyPcVWG12/VxT+SPgTRcf53nsxubLt1oG8S
HzaczWkt4nui5aavYz/Rt6yzNQ14PI/JgfTiixREbxzlJdw3DBf9XqMMdfWqgzGK
VbWVbNW6ZNk90xH07FyDlUGIuwRBugTbJD4EBVuY8o0Z3CrriGWa/DPygQGpfO9x
NSWRM8sxSsfH16iRYgI3/J6aofCV+SSxKmy6fdBZ1fA16bZWH173Z44t1Gz7IVv1
YnGpvggHY4ymKzg2V5QmqEIGre2lDL6bJdn6d1SekNjBfDV0dKUqQH3YCDuGu4c7
D5uwB63ZLC0rWy+GL7hqmrxQyXvnObbUanajf4e9lbjQtPKYemtnbsGPv1kEPDM6
MISrCOeuw40EMsnfyg1frL2gKjoelrgDAu1y1Fla/PClmktbH2gmq393gq3NcCai
FEFOm06qtk4CIDyBBpCC+WmzeTNdUurzohZhRtAPRkf/3IQlNeHy956oq1qz04Om
szLc8DgYWzi/OB+TEpqBAD0cHB1pTPxoat+ES2ateh5FREG54v/426CD4Qi8ME6U
LmtZVlXvBGX23NzD3UNcxmPGbmSsb3bSu5m+nWeJICh3VSkPu9KNBTmN/A26oKpz
CkMlWNBrng0qYF1Aqw5DrvZmAOTQ4AzsmpK9YYYHfYI1eBcc+pNbx1YmkayaJ8Ub
q3AKaEnARLxGq+XbV5UterHBHf++G/+BbBEmt5fngiC1iMhGXXhaZN5FtSyLgV+U
7Rx7kVE1h8Aemjf1TG1+ey5dC1J0b0lLx7Ja/UR14KvkuyjCxERPIeJoDE8/1CBH
mjrS23NQ71gCOQ14tJ75/adFt5RbBRG6JTbiHMVdveOSOyFenKw57+Z7QVQSn54M
SXN6ouU1zdGYz2UxJfWhmdNycToy0/YqwMKqa158aHdTgZepX4otCWuLlMxGoNTI
TJgQOeBdarlP3ZGTP9TCqoLWfGCMQUzt+yvl3xkOv9xzHV0DqTrtQcChJQtDv1f5
jIN6AMbQ2noJfOeEolTbcuh3paIDHv3ed+/1r5Z3aw33NaosRc0sMJtGIJcm797X
6nk7m+dufXzaaizmsbyzpvCidB/Ju5Ykq9rY8Dtb7cDwsLMRTiR27SLcSNC/+l2t
GzQNi6wWtcY/wEyfgmiMMei+WRd/mWUlylo0seiheOv3nef6DrgaLzHVUF2mHGGW
/zOvrxKgcn0oalqNs5RFJH6zewt1OKC7pCY9Q0eVVTSSFTaJ8oFHwSjC9cN9kfGQ
kV/TSVYH0NFLA+asWrlwoAIGkbIRc3PIoo+G7/iw9HojmsiIrG3PbbAoTKTugUYQ
s0M9QRNNyrEVrefKy2OeLaEWQ1gmltATM9lVYEDG9BiCUUgGoyDxTaNzu687zgxR
o+wi5t1ia+6tCHnS0QaAybjdhQqdSHWBDFOW2MG1Rn/NKkwk01bC7I3t6DK3JhPV
ukX5SJIrrCj3/0i+N8LPOARFC7VcFynQhBKBMOiOPRN3uwj9wwOILNwjMfv/yOBa
egqZyA0BTmjcB2cJ/uGx0vTXJW29DB7++WMKofgOPiCDsoUIj10OYH0+oVOhqEcX
wexrZP8b/RI/cGeXtsdumm73OwgT3zEUdZOGtYlzdNm3I+LBYU005/iSVTW39Ltm
pk/ojrRsk1CaTlfqJ9Y7CFwrYql7azq7HSjaHQ9p0IyfET2HjrvOV0OeJjPWX6oN
UnfwrqnfL/m+qpoJqHdyK/hKyHlpQyiNOSMF1+8m77SqDHpqF2KqThkmcokshmXS
Q6QMRrMYvJkw/mGu0H3H5NJQnKmjmOgD9iNPQdbFiwIK2BJQ8kqHdvHhA1DrKVTC
SNh9v4OqvqNmUy9BpdD6sQS43ljLYQelt38wvFVJgR1kAuqeAsLzZBhMVCHyrBx3
WWulMnX5qBhQdBQtq95voUrB1mw4+6P4rWDDpbakJtn+R3qH7hMIXPXads1Ijv1E
PWAfVychWwtIrtqKZTVKe8n7x69Si5aAKg56K0Yq3zZlglXDDCBdRQ1lWlp+XrRY
fHbrhCTkIRDuE8CMdRGTdIcmDPBn3a7vyuGsw2cCloq6kzBXyobKNZi3vqxeIxSq
bDYzuze/o6ryBM44n/n2d8n6Oys7co8bP+o0AU1yRTIQk+qxWws0gyFAE4SrgBSO
Re42ecKDSAG/lD3c01Hxi6RKApo2KHfu3njCZr/elAYgpC1/xGafj28d8RvT/g0A
YvbMRtzVOaalmjyWE0KCMZ0AFgGkMv4X71L08vq0L2Usr5FznhWp/dL2fRVPtLpd
pAx8W+Vyp1fzSDavOYPTrGaEh/vzVoTmrPifkwLdoPS3HkHnPF60eOrfnsC6oGzb
mEgd8uGBZL3xq/VoOueg5AEAgR3fFkDU1p03JFR2a796X9Tlij1BB5Mv4LENgpyX
URVTcJi7SH0G/y9G1M9UXNMynPA5vSbmuf7YPDPNLjZEsI2QOu67dzz0YNGWFNEd
Vh8+5lJJXQdCSR56tv9E9w54MJBGz5mgBNRRpGEV9lciiYBLK/zN4ChlzjPzlARZ
Q1PEdfWjeVF2cP0C/MJjeZFqpF9SPrqCxcOp4LgCErwMtThyJl+QCaSo69qe/VMn
3b4/tm8Awx8CYBCt7HzWV9EJM1yjP9+b7BNj2PiqphgKbF2Sl5Z5XVm1G87P6PHN
AKQFAK64Y/AUGN7IddqaqPtMNNDY2DZxFldPJVQFqDYT+l+8wu9dRLOBjaDvanYg
OhV/aa69q281QctHGd92t1QI1ZajuE65v91kwbO66rGsOUvj3zvLngTXzeYUyUhq
ruEhzK4d5v8T4LfcGvcPqvZUkW52yJtcJA8CdFKvsw9XPo7lwahRxIKAE4EFexC9
oF/AgIHlWJDh7FHsV4uz6+BaUJhk9kCcXIdqCpQCN+sj7W967XmhjH4LGKeRgJvn
RL7ou9mr6ALETxCApxyfJR0XKAgKGYlB4glU0AcNe48S2JK5z3NaLRp2paDlFRYV
FUrjupOntuPzkN1uZ4HGSBzzhIeZw68oy1NApmTsrDQ4EVm/6Lj9+CumZdF8X70c
RPddVUUMIFQRm3AXNKxnRSP1P5cfw8YIBIdOJNv/4pceHdRXVO5hdS4/6m56aYd5
VwD7trdapWkPol1wNZNzHtRMIcToLe54HHy1m25Ep7WgJOwLurWDI+TaSCvfS4UV
yhsZRYlL4KlF0UBk6SCET0xeJeAALCbJHn1+vRlkxzrC8kAGddgSPEfVSfPY9+8Z
jukM0WybCc+YdP0p9Jg4m13Td3GknuHj4f7naNqgfu0/rz8j4x7Ko1PG9NBiYjfp
V8yCUeeR6oYTdgrFUZImCd/uWIanqpw2auYzQfsFsuBAVtPPvd3FvZ92ZsJr7V2Y
crysagzB67WsdJgXn7B6z9RdxQ2JgAF4WR1W3rSzm5lgBLoWyW7YtPnKEFnLnYF1
YWl9u8XIZOaxpmO5dYu2aVC3FN6A9mFEBXCIJ5TiPhRaikpGpIc5WPQ7bxhc+zJf
+UwRNVUJWbeHIZgOsOuKWxmQBEVmVgDbhIK5k5b9oZCCBbeHBaI7U2R8qd6mDZnH
ZnGWthFfqR6dHJD2Sx/dD7Pvdn0APr5kFKH8kYgMf8mxHe/PwJXnuKhilUh376p0
oxBtlEtAZdcd39eez3oa7xHhGvu9Fn7CZbOEynZKyUcq2jGWvTsrm31FsEWYcccc
woUVV7syDMFWDWCvo5fGImeOfzeXFTLhimj9fK+wfGAziIGrqwHpWMWca+dEToUh
EveqVVAzea/Hx3+h8JTWfjzHZTMmKduMw5M6BM5AmuBDO9zr+5ZAVoVBkc9YLraz
EUsYhFfzuHZIuXQuElnf9PPf0g3PGub9wcQsen0qziWVaVNTxOCcXeL5kP4aPIpS
gqTT7/KH7hdQHYQ81jWv6YM8z72K+k57Y1/uv8yTwKHygmiCYACRTQ2rnLfWZInh
qN4g2SRTMFDr95zoefzANcxAk+8j3u2auN2qbbNNJyYFxCb8xf3vLSq8h2imp6k/
DR8mKrA0yql1asVhIrQHQ2scx146YwSd2ofedQl8A+obyOLohASSBVnPNXLh9BrH
JHfz0SSQZPwDQ+Vr+BZXg1OW4HOUI97+WQfo4INJNzMDMnC1uco4kkEdzklKT+vb
oRDRAPbf2St72vg3RoT/iN+z/UajOkeUVillk/MaKKaGWy9hpbVo4WqSTDY/uqcQ
kLmoh8FvbnWazPv5My0Xp2EsRYlF56WjfjKmV4de6zYfvU/JNwyGe3TrmmzecoxK
ZJapQyoROkPPV5CcRLo9/NxysMA0YJxKpRnLflzfXJJ6OkoRNJVXkNlEHuvGUKG7
0m1AO7watWF0AKCOQBrb56aWFZZRc3KG9nG5glwRqR/8b2UOR4+0grmi8qGxNGTg
vqIfNcjzvqCMB2ruE14V2QnyyGi60aHzu+E0NyH8lnpW5ALXHZxIwi5QjSjCwI19
1SgB1xpySnOCSXK0wXwK4v29OIDmfF15LeRgosuBqHuYKoZyaqk0piLKlxp06q43
V7vFzalBcn09fX/iXcT0wNMeHZSoB0ffsW74/vLwL+xMeXYLBEuwWQa/QaTCRyHO
rU2rP+S2p+QCI+vHQym192g36qV8g0fa12FqF0It3JPtdUvamB97VQeMu0cpKhYU
yY4vh3/Sk5PBJnfseXcWZoP7do1jPqhDcPx6hJeqOp5bujEq//b7QiQXSX9emT5g
R/NUtY7+ixjNGo9gz+W25ForG3gF6NKao+XMr4aLsRodzGJOSsun+2I7JsA3qBQn
legMlhEqF+pUUB3Y6w0VNboulX4GrAvdfRU4qk6g6IcKzYB9OqvhSlt45Kp0LvuO
nl4pftCOHHmPMkv4Y8UKvqVthGVT4nb0z57U1dqA8XrRCEPcG4jJMc9Jdszuus5S
PnwnEVOPs+yEatLwLESVNIkEu9JiehzLZS5e8jnzeRGdphZUVsdPNEZHM8/2THHI
nfLfeqCyafpM4MqvZWq0vd+TQBWNORxLpZlE5cnFZPUxpBu/m0CIBFV9Se4rZF+G
6JcMKCrSl7F7NIBcL6Vbh7uSTUedJNu4Y0VlCS45WJyC1wHj3xgXkXdY7VblPwwN
Z2O4Mf/ectMKUiu9XIsGjNL1pTmTACA6XzzQnTWktbNTzNbH5LNlr5HQZyz0CFOA
VuLRwZv2QOarW+VcPtHSLdNqTUuKnywZtvTs0ReQuPTjmcc0BHBGsUvDvWBuoHQ3
XVNq6kC1G8HaRkdGpGS6fuXpdqIOjEtkZIIejH8mhrJHSLg6xNet0n/PzngnQQDd
u0XbMabkZIXPA0bkKoxjaXF77WNvU1W7OF35VOBkd6+2r/r1sYjXZ4oR0arJXvb8
S8Dgdg6bKqODMTdAyFyJ+Al87XgkTZUpkr8wP2+LsE8aYKfW7CrNuJAgV8UXYG1E
sj/92iaQO6k5jdQJ2CkOToC10uCLAMcegKr2Tl7ElO3VYthC6wmghole3z/neyME
nF7nXVmBn8laGA6pO7lniwwmA/1Unjo0gvtTJ0l+NcBo4vcZNFd7+UepX2k9ej9W
tQ5mWF02/3qZ3RseoXqxeoA2e5xi/eZkK3dcpJSpgggV9+mF8idqFE7BHBNB7Zqt
tahDZG/ydvtunBtyXnaooQCceVifMbOuamxiT1sevkI5IbBx5lTMQP/9TJHYthO4
7bgch7+PMP6xJ22aDQ8dNHa2LXRa3RHoZ7HpbK4RCRUV/8ie80Eu0ybpPIvi+IM6
aQFFrkMc8VVd4WsezbOKVucVffYhO3fGafhgQBFSm7dW1DnuY9+Kl0bxxQy+CeXB
a8Vyg6yFf3PTesfdPmER8WoEWxvzYsJHwls+ss0sEbsm3ku3pfCdnggCUKEWDdE9
LGHVzjyyNhrTcWjjF7L+bj2mPEYtvMLy9QCJLvQEQL7mq1dZJXAuEsKPMzih4oyv
oTKlSb2J7dW6xUoExp02LEEpQn0nfTLsTm99FdwIarjo4eVc2E2GehUwpabHxrRm
ZnTWTIqa0pwCM1XraRqxiphGgIR8jc2UaY4TlJfAvvxo5tQfRtXma/5IigKWw3YZ
TlluR5XsuAF4mElr2TABrfZFW7qILjul8pkC+zGHGQizdcSc+eW1jVDHOIxFaplx
4QhEEynCGGOL9kZ/DBCsFR5CcDxKpl2h92jy/x6mNe3Am755fa97iM0PFhYQTpy7
eO2o7/ySe6ChN3PnbQ8WgYju/bubMSF2dJtF+Wdq4Olm2nys+6pn1WzIvYzkK9L4
tOyikSaqFWS7owreiybqvVDaWVXqy9dcfu1qRkFa3xDsJuF9WgtyPBeCQlHh3Ej2
inoX/1s2qAIwUL2S6p/trFxJh22O4dSPUoOwmwZTLX9uxHsKtdrNVBttxc3+dSyT
/9SduVTF+sj4N/2NWe1+TP3mJVY87966m1rRqmk6edtAOJLD+T/5TKCChE6ml88H
KCb9ImaUzzln6sMOTzSZZY8k/aoxTKvq9V7LIAICqVO4F3FehkNhA6CuFpr9LvGY
J2fnRjpiDIzj9j4qalup1RpAS4LaRMhEAquTVkOIae2z1kU5xkLMz80cfTRYMjDi
+06RABQESrsL7Z4uEaUemzubpZg0ODyyCAV9XR6dK49yZEhASU3DEU2wnHABesEG
1sZuncYQ3xicQ3CcaqqAMtSv7/AKUzSW4znxf3ewGsgHYTI9LvpDOdOCNDI+Gyy9
n6YhjfJnR+6sD5tQzit+bX5x0l8tcHyo7+Fhhx31USQVvnBf+g2xsTl5WrZd/Gox
Xf/cWT06ypWC5Egw/ny9kiEKdc8+if2RtbtcUSWpbeUY5ValzJaApZIqR3o2WKeG
4nFHdoRJ6SBvgzEYkHrqZmrUH4spr9iwBQB4MehqUGDW1l6X0zRjDgAAjZIvMBi0
p7a1Zb1OAS2vFM4+ucwsufHlK7xx6dJ5oKGKP6PQhvv94Y9Ciu6jPI8VBnkuECFr
342gAXCxdDYc5lAIHPS3/irrI7TAQDwn3RSIAZuiUEiv+0MqQm8FHEXnKWKrKk1q
0T169HI5kbbDJCU9e46fk3AvwlDY70M7mKgdNdnGP9XtToReXRzPl2pt534jSVNk
2tm5qQnDqouhmUzuEptcNyy+2mkIx4kh1qsbqk7inevoNZK9kH1UxcifsgxnXXRC
dU5vHkrL+t+7pXO0woLY8UN7BZ0b8nEgnFNiSYaEuTAw5UgdH5stt4R5Cmtiuo0u
IHgSZbXCBP4IEk4yZ52r9PvtApepGf4qCIGkITxoulz+cdUi3rTXdjo0CTf7m+OI
w6h1kj8Hhedhlthcp3O2o4OBY6pL+1EwJQqRRPD4L6ovDFiuQ+V0XvFR9Lcmjy1p
olVISV179vNR5igN3IqnXTe6IzqGBIMx39Zsfs5D+M5FNuXYdV19/fYc2FVn9VPQ
b58AzerXCF1nZJxGWhLTNKojJEyLESe5PEni3tPeqwi/TmKe3OjkBXnwACcjC/d6
BUy1Q8JEQYjGjPCBSqh8tDr3j7mlWXdu9KjO9yeJBRpZSKZv34ckNobbM8rRGQ3R
z/Fn6bJXnOXXrmySUQwCK9clYdXTwp6GiZMRhpIkx3D879mpcQnAX0ouEAPrTMZ4
rT13odniXMG+7kaHCte64ox7F5Gds4LFH/5P4Qhf/MIamtX7oSO49vh6vdguiHGt
qgNPSa523J/KWk+TBTLVw+tg79cVhQmn1sQswOHjZSVL9UOtxJ+qY9O3v24J+kg5
WW2gQntaxIBovSN8mreCIIp8hbN57axaPqBbfD8Vu2VwBg0/496zQFKHA+EKbKB6
1ARuFSFxWmXGP9OkNA/XzIwPVY0GuIPqBTfqPIINm7GZCuu2jbPP4CXLAsIi+u1e
+ebkwUgD2c/Q0KPfOSgJucH5pCew8XYnGaj2/buTpwB+bjYd/mvPsNzHlprmEw5L
z3UVDme6RvarYvLNKD/p0mQstBeCYI/1/1UVUE+3ja3BmwJ1rOFLpXFdLaou7ADL
NOzdxG+d1YP8FkZaziSXDABuVCIgWpbJAgvuq8i14T9PKIVJ7huaZhXeTzQ6QBY8
aMbEA3eM2KLUHUO2BgJp+k28cWj+nxktE38+G1FiHwB5Yyc3P9ItGwZEdRbTwf1R
ZP2s1QgBwJgjw0HV3MtLA+31C4SYX2/kqdKvfbpfbts76lKC3rgYYVOmTrva/Mmj
QSQR7CTECxjYYq+nku9/Jfg3kYjNnX6DwMKn+vsmxwwXuBqCuq3OcTBnk5JHwxK2
ANLCFDEFCY/E8hPKfkAAu9iYxs939xyNk74zhXgqFENMx6EZ4nShcjMb2SPjfinS
xK0IgvXOqipfbm2t7GgKi2rd1ZMfqXPii+gzliYIPQTvL4X7UzjWiF9/xQCUlldF
Xtvpdgo7Uuo+xDfN97dIkdLxcQWUDes3MZvHcWI2uYWsm0xIrPSpPM80/Ut2xhHZ
VPFc4gvqBrOdKsB8MoNHLGj08A9grtE14IjGGndvQogrs4STsqoFnN2rFDrzkj3o
XRi6l+EqNcb6TnJf4qusbU2c2KifW6xJkQ90Rx931l4ffvPyK+k2geLeYRjeVaj1
EfYjf7oDXFQyhX/zTrkhpqyFfwtGpetb3l+WH6eHhuJMPOZKXth5zdeWJw2AnjmB
YNaVInT3/lNzKfJV3DWMhvAlz2WvLSK2sZ+QQQIcO1EeTgRx5k45qOK3FF+K4SdP
8VmO5bwnz68QxDqKoOD/zD56XOYnt+GyOOaJg5AGUMjNQfu39aBR3TTN628KOJeU
COc66ezeSY3gHBwx7DZpdk9OhLM9oy//UOHoVQnE5dd0/L9DQYLwbOMcqHqNT0wb
9DYxRa/REbsH4V9X6E+eJiEALui+rXALRqA4wS1jc8FqK/7L4CdCLR8HsdiGVGsg
nRckHItdmaa3Ua/OUQ5h8TXnId7QA1uLDc1PP+cnsYK+g6yFU71umfX+voonqQ+5
IEDzizIWgpNFJuW1Yu9i2Cw9x+LJjU07Hvjoj4wwBWmVBkqT8eUVhXGYxJzu/mQC
WrUbkICGNOdE4IQBIlfT68PP4qA0GhOhht1xHocK2r9x77TP08O+NkA3IaHCsByw
WML5qhcB/eSTN+Hb0SXs8puItZiaTig14JDvYdy1OfFLD06bFvsmx3R5boCj3PrZ
7ZOnLSnSK8zxi951bcbCxziNMHC9kGCyxVUeNpzX5R2ncB0YBtEN5k0VNjJ0thCT
8N6fLo58sqWRb2yV0aveHt6U4hKtFfwJeAbPmfv583cFB8y7/5HahcJ6u2xp+9Wt
VtoiNlqVzbFx6SPiYugRg5TvXm6KfQJkbwY7htCqG0wNNGJTjBlDBxUqAyhIU/vm
4p+QYcmfNSYK3Ci9RrDbSPb0w80jvi3z7vHwj6+M21M8pQQLGC2yQM2ZeaLkEbt5
guU1A7QuN2Smm1Anv/1TQc+cseOrPH4hAglx5IjXiSQWL69HPTbPWSOVr6+Kd2az
rZtJD9FbYtTJ9nrtpZl44pMi8mYDo2o++osAZ4zzMuWbu59P0dATNX+/ftSiaZst
vAe2BMUcxlHCdLCMmO8LKo3wI62+2xhCbdVTw6B1WPZSNmH5rDV4yaeX5JDF78dx
xbozzLyDK16QEKlCYDORU/rk1k9gGJ8h5BradW7JuPVBAhCpXtE5YKQELTN0keSl
aSuyr9Sh1Was+GWUEPdsRIy61CIG0byOu24PvL7FDCWi4l5NNQJpYEhGWK6P/1LT
qoGuyX4Stx5PGo7a44O8f2OKbQkqSGGzeDRR1y2FUrcobxhhont5C2vnbKNM8RZE
VbGqzvho7Me1WtkIyONl/E8TcYYWRcAcZs2E2vqrz+iCws9catprqUTSKCBT/ose
5xPO/u2raRyynNuTHxTTFMP815KAValMZsZePoLR1+z7x5K3yGRTYo8oop8CTlqW
SGdqP50WW/T8FsJHDuo/LZd3hs5BOROMl51DBWY3zJ0GMgjksNbnaiTYs3MMYCiw
8aNEBWqIaI919wdebN2DcztsvGqe72yKFc3IjamSulPYrKm0MDHl/RfVFCoim9pE
arqCDeSzq/dN1j/Erm2gYdg+zbjnoticJWTGHaaPihdvSOV8HabkqQIWfOG70mIi
iM/3Zn4PwcNqgg0mW68semh/NsdKTRhfSzZ/Sx5k1PDkOHV9ZyOKCukehWF3SIFu
rEWcMLh1FpsJXlCIkOjSvlL5ileX6W3/O/n2ND1z87mtvr4b3F9qFKlL0HvGOaW4
Cvu4Q+Fn7oD/WThv6xbaRP79l7FUsdbwyDKGzO5H/KsPD40okVnWcXUqz7zhEfeh
oQeIUcFIShVmtq0e9v6cb3aqwU56V0aPt7E+8kmxdquspkbl0JlCyHn6kUyobh3t
NOnqDV/lfRxBdVgSOluZ8OAvAvmg0RKBbdn5UGz1pMTCxViJzlzfFCVu5Psd5ZOJ
v6uHHjqMTMOvPFM66N3pspCQjg6o3WDLybLPxcfAyujtqNg+SIOOeAYVraV2GPqP
YS+T7c3H6RKLD6KzSb7c55GkQYL+yfKa0euhBCHpD1ZfWUxaouWenyjtUxH+FUh+
FpC8w9rlz5wQcDHKCS9rgyfU6eIGvpn+uRlhyJWfd6BoBBDtNjYyeq2fHZPCzrYt
lKVOvqKXF13PKKOZLXzqVs1kZfmulH4v2ZRX7mSrXZld6G+CLqmW0XSKZvE5Meib
qLprbGmKqyHR4HkHG5NExsoFGQaWxfTaoPZQ5RaVJ/3oKAculGdYP2rsbKk5o7vh
szAVpq/a/v4XMsY1woJw0V93+Nf7PY6cqtzb7uF4a3Jo1bq/qh8IqGm+7pQAn7Le
nJaNoJggfk0SKHDOMM0KDsJpVp5ReVf+9NspN3tv/ewg/E8jmf5z8n+4gqKI+7Rs
ZjRWhyDS0x4evbvssPJiZZ3emD6o2b9sU6fW+KpcC/XnzZeQnugcj6Ev22CRvXrB
YwytZh3DLrV0+q8C01eopAL5VCME3ej9sSykZKx7oLZG2G5NJ8Eps20o310ksvkk
2CQ8nz/Q30tvZTTG3huA7TQuWEFsBDJR7rH7Be48KMVBMGGBVgraX5shqbvo//0m
0ODggfCwUixSow+T/Z8h4/lLMmZksvdaBKKrx7oHvGKiOan9kjxmBaR0JY/r/FtE
H0+RTPczrPv6CbozcbPBH+Ovkyqnq8gqJ9nxV1Un+1/oFaHyjrLvV1pxdqMscajJ
JjhN5Sf0G3cioT81gJ3TMniGYlOI3jv23m23K8u7fPrFgYoZA/UNL6oEdvk3Unjy
S+t757svv+C80mCu0TtAbRSsaXGEBWDqAF0GU6E/Dx6fH4K1Al2gsZBqzHL1C45I
siFhOXaNosPFZ/JNMhsSfNTwmBV0heE2pmnXpD59+HreRxobv6q1g/4HF9GQJosZ
rXQMA61i4k8icUiZnHC17KLIwiO1aohqQ0QXGPOOh0XMefa0O9JwOwZvL5xHI9Ka
8anzj/gmhs9POqrFeDY6Eg==
`pragma protect end_protected
