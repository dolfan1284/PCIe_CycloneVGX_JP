// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hz+uHTXWmYiNHo3+htThv6/kSZNS49e3LTnqGd/I4v8GA1m9ZUwPqQ3GWfIvdckG
iXXD8BeX7NAHQlUJagSF5QtG7hAzmeO1IV96w3QgehIGlGjcEtVgWk7pjsKr20U/
YKKRVxRPCsgmxKp6+D+41OM1PJ7SzxHlRxnkj01Nos0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4848)
gPFTZO2/P6bBPUrNBiQRBI1cOxaHuVWdz7GBnQIpw9MZR6IPWoMFaYLexLXo8Y2c
NOk+Qkyu0FX2DCCrqAj++GRnV9PcCylaT95/rffQbKINsOfz6OZByJXLy1tFJQhT
VNyZ4CxD++DgAavgHuZ6i4YzTeOx7FUfhtKdJm8tvuouwazfPkWVUDGgVZ6JYx0A
jYRtde0ML4syA9m5lzTzFeEYC2ktFf+f+oznlFzDRG4j/C4umuVjpgbRwptl+uVz
X99370qExeU0We2wePk594qtzDGnsr7+eao+XmCd4IYXlkrH3l9IaN4jZN7M5D81
SPQMP+4SjS5kmHjbyHOLy265sHYZUEGmen3EesOXC+xzPq3Kfu5/eOv46Wn63YkL
XNR7xZbhcvzrTE8qhFk9t/4ING4sJbXLQMtjDL/tnw9yWFWNyTUROgDRuesD5aaV
A+elJfuH6nESyxYCTNNC10vO+He7SlHqqKtLnfT6J0pwP2uYfxpR0BgMcymtiksR
N6gqv95tIOB/TNdlkLkbpgOfKYeZKcgYLNRWn/aS+Q86GOI+q7Dg1VoUsGSIcUj2
yEsNSJyFya/7cfGW2qICD1O4eXRdpcjrOH6vBWagNvjniUH7HmultUNqmfPaNSer
jMZT8pH1tCrVbekMazUW206rV3zxJ5bW6G2sDpjKxXjmaRUurNmYOzqaAaXXsQnB
BUHAKNs+/w302whk/ox4jVZVbAmfOL44VMlWICMP+hpcUp6QVAD6Nm3r3J72XCo1
inh0oX3Fh/ocMeunjprmqIjx00SLkNyX+6g4BNhhJ0zkbYrg7QCAMeE/VRP1MV+T
c6c5qwWGJQXccw4MJbL+O/ftTOxgSseGh6K6UVSa5yTS6spUcz6g8o21FkXd/Acc
ldXHQCkWQLi6w0R6OX0ySxPbKq8Twp26aG5NM90IbjGRYNDHQ46ChACaDRxZewdj
ybmSQdgIiEyqq2PxmqX3Zss5nP28hgGHs8AIMFOuU/gT27L1DbRGV8s66t7qIHBM
Y5OqNewXEtPUErhS2Uw8chxrjnltwdAwPCtkBsQOx3xSfgYsN89uKnY9vAIYBWgW
JGb8vm586C7FunvEZ9hxk5v3IMm3sZqCnGxxI2CQVv187UAwoDIF5Czzt9nIsiR5
mnyqTzN8+sQLDAMJtRBN3eOJER9vAq9w9tiLq7J1Gk9zFNDenA/IVMnIeBDlsrkc
4YI4uSOTWPUoWh66elr8P5vzG/C5Eo4laFDuy1D03YzwFtTzWmV3R50GK/+IqkxN
5+K3JWXTy2mD7qV9/h4nMIspoI7x9DTG8WO6u3rHwVvRWHQc6P9FY8DwnCDjb9jV
a/N6+Scy/YQ0pbEpK5kSuI8Jbt2ybOaKXCjH5bufo4G/qDLhbCdZV9pnOQ8oRkm5
1Z7bSwLf2Zz7w5Bu9fjMV6x+8BF169SUoGNHXRWa+hpM7f+CjnDOliQQ/9SFoYzY
ZbQH7ZDwtqOMTDQlOtuwc2Nb6CsEr+TIidocQ+QjpXkXTHOyGIY86uu2R7qpHtkO
8USPkbGRi5aNVh4pN8u1c/xTu5Ts7FIRUnfOvfJ0XINF8mf+mbwjLDWK7+zyTcRc
NfVENzreFtbNL8xoQ7fyV19q/GL95YPo+K5PbwmYnDxGGq/Cx904CkHRyPY1xEUn
95eZxz9vHveeT8+QBuxjaro5rpbKsNp/AY8B5X1ms3W7CM9whEx0BUEKtNoyUJ2R
Stdgdn6MwZzVTIQIGgJCHNTrlrKHi9OUQN5Y394pDU3ws52pFcFlieTRSQ/r7kca
/NwoRYeIEuiGZap9jfYWHpNiYszPmEL3rZnqtN0ztSoy3cNa2iCgo4Gh2jKX5yia
M4GisI6i4Q/3wGO4BSZzDOO6h45YbF6PpdFnaQd2o9e8N/p4XgCQkafl/vgu/GyE
FAL20GZxt1caO28/OqMt/bcjpzdN0+Hv93A7RGEVEgixCX6mcUDs8YBUssfj6O1F
/zBQNpi7G6xVZSkZ78aaHkZsfprG7A+Fae4W55BVQxO9G6LRGMZRkVbkl/TadXaX
UKMyBTM5OBCMkiTmVGE7XH1IRIwi8JmrrNDNwweWIE93H766rRxfrxcB56+l4GlA
AbvixeqGhNvIv6J7PYXtddon8fTpuWbpws7Tqk3I9Eywsggic/yIUYmgUtE928Om
IX5+LyceKgZU4qZXFqLEx0TP2z3H7w3UsZ2Bd8gzDynGiFKl7WJ+rQO1IeZ7c+ZF
G9rlfrM+S1CGEZ1I6Pq1d6KkH5GrsCkI1zf4TljITpfdQ5E7Lc0cokbWQ+1ULjDb
k1YEAl4ER4u2uBGob+YmRIdm/jMK2i2Xu8RuVtTc7Qg6gcTZPQvZ5KnmCCLbaEUo
CX6jcSOKry8xXXdAx4yubz0IY1OdErMs3wYUsMoy8C3JYB2QpWvvnkhm8hR5SnFK
uLFhAhyqShFct+CmCnrPGepECjOwVrRD9/ZspsP6m0o0/Qn7pBRVp1mnCHoaEo86
RgGMwKVBQbnqjyYIPogVzFR3yKXpphUDMQDULYf6lC/slUvhVwC3C2z7vTAVwek1
vAOobmQXwTeZESdRWLg5nJCT4NkOOD6Y7fSg4qcLjUNNr2bymGELQEjGElLO0kl1
/OxbBJFEVrQVd/zdS3DlIvLKOrYNNeY1sotncQF7iq386hBxZYCHOamiYgW79BSL
b54o0kmlyV/0E0lD4o6mk6mymLxPp6Eqa00e6iNyBRPoqjj3nIEtVLYzwwdhn2Ae
WGActvty0IjxcUaVveSt5tMRvqX076O4uawO6xdC6pQacsw4Yb53KciyyuCOehzO
ExEa4o52OG2aH/Z83fU1Ot+n+bObKTVbRc1AcR0obf6J+xNub4/z8O7kMAdjx9Or
4rY470RVmh8syBALyNNAtUdq7BnSbuzX/MIJc8iQs9xK0BKWhS/DDSQyXo75Y43B
I5Ch+AvFVrZyTFZ+pmGtvuUDdvbfs1f6VHiw97Y1xQU2P99LVUZVgV9NzWtzt/in
GGKROY1H4ig0d6DZD5n6E7dis0P2wgqU5vHKK6Xl8PTtbtdoChSqDvrtxxIrrbgs
uMvInEP5t78F/dXlbhq2dZZeD7udH5ggzhn6AVIqyQxfswcxdnkJ5hjQtWNcobXB
Qym94wS5CObG2QwElIB03KpEvNsz+88Q+63x7c/ZRg/8znl+2loBYUOoZzfthXqL
Mknl1SS5DxuY8B83GXKuq8lO4rc8DbWf+2aB1DxQOaW0NOUGLQLeSq6Zveoo5/0R
30AmJefd1p6+1YiB/LXU21YhtcdsgLUJTGCXSU8LKo2RJy7LEH4TBMYzW+wC1m5m
iNiXJZ/bG1mhayPi1EfyUcUgxB26P+RhMYBOQYPMBsryDeHY7iAzwjZNaNgLUHYZ
GGIkuUoWGlA9AN9qkWsmH6HMwKO/zSoz5uZZr+eGWlJIdmdS+fiD5i9+O+h8/oKp
hPonpJzKXPixpx3j+VQRg2re/Bt5V3YXczonqY//pbefUCHM+zuuLC96i/HADnV5
CamZvTgvcHAk7kLPfSfAisPw+1ztgFPBdrKJARkYjwbqWpkfEKCSF3KH1fca6PWz
nv5YBXRxW3gncvCwf03LvcQC11q+XY+/ejKZX3+8xhwJ4WgpX6qnbZy+9aLtAWW8
dZhF5KW3kTkzCJuhnSDBBVl+AiE84Z2K8d9DB7EpwjQlSXwUNjAIcB8SZrQ9TITO
jReupjP03qj9I+g2Z2gbTRfsDmd88VPE4gamICoKLkeeTSxg73r32f3fkc7ts25w
kRgM/cYQhePwxMK2epIacbXXFM+2DpL2lC203Or2NZ/dHWem6ERgeA5wsWOgM9bX
YH1Al3aNQF5rUpnPj48Sc4JjhIJvYC/WHHHOUViDXPX94zvWViT7h8kh37GdCDp5
yL/PdtyMoSCa0cjnh+wrzPxIGkaeZnnKamabVe1G2/4EDyWeFIl9YiEHs4TPD5hI
rD6K8HRTWGhnyqoZZg6qnjITkUFWVi/iC+ao5kII+uVnjiJ+qNwNAqxMg4AheWC7
cBiOl1eHr4dO8c727NqTIR3V5KDn7ngqK92ZNmv2T/u8+YXVGhj8Jau61WtYztlD
9mCBN6cXFXH2G2cle0JAOd6amxN5Y6imHi9HNTt1QQB3fBN1vBYE2VqPFlaKgAYx
Edex+sVvs3T4hbfJnGaG+CjdRO9gOqPufmJMPjsNTiBtBjLexTLK/5BAvQuO/z8h
9Zkisq5lduQauTkGgkcxa7nBKDSmjAkbsgGGgQuHlU28PIolUZW1hyYEqZFQDqp7
16XNIkKzVkMq/5RPJUeq9UmAV3pGKo8fzBV5L2oo17qnRYIqhZHJinfNtO5i1Xks
WD2eRCbfysri8o2iCbKRIwjPnAdYThRpkkYxr7223IzSTgQlRkH6pIi96oqBZciM
YpQAtX3BqZHfecLN955vdblQkGY4dgI7ovHmuq/vxkT31wvXhTAJEO3hCMdleRfR
0l+8hFIXyplbmhktt4uj0uDvtK/S7qCr/h9nyXICfXLBQG5k9apCQdkxOFailR9U
YtOghivQP6GTcvUeJa8E5nw649zK2niqDA+LZsKcrKXA40l2pruc8ZxCI9AH3QGW
R2+mSQgIVSf084PoDIEcyIUltQlre9JKvf7lDBbCi2NQClfz05026F7ONE4OKR27
mF2ZL5kBdKlhU6XrXHV+WmhB4XhtStWmcdviFtAzCpiJjSjhSgm8E7q55tFYTedn
KTrMQTjh21Q6u/CJDVQQrGIbd3k0tuWoz/vfQ6iMXvwvKxKFxSjRAnzp8TGLyvrV
vYhVvmOm7TRnGfq19I5QUscuCPvgquUQz4rTgyIztWf8A/diMnAb2Wd6LWpHSImw
TO4+b2AyPnK5SMIAC+H9AZEj96n5TRtsgslqXYcCyff5tUSFijDwR9CeT6O9I5Wj
G6mns2wU6emPCemReiRUIPQkPg0iCD9mEORvHocIe2N65HXSLhrIQ7/Q1+sDEGa9
MK3uFBjnLfbasXghA79pY6UW6+j7heyPS4igKZCInlp+Ftkra3XOlikGwE6YWYM/
vXh3EErt+3+qTH10oWrNK7i2tS1AQuSFGa0uD5Agv2gR4CKm7JTknVPQd0/uttSR
nyMEGpNMr+EUS5nCCT6dcmsepUijShE0Xu9FLWlUAGvPacXD9zyJzZL3uavQ0n6p
LU15D1gR7LtVzGcj4yFvcUjtJDsZBE8Dh5OzKlfNI+JBS/9u3C+rlog3uDT1Xpns
BwEC86UBuRrYFT9B2nUfNWClZ5pK0UnNJZVL0ILPh+wqCAhVNJ+ydix+56UIIQ3c
s9QlPZ8aMxrGIuF/bnRK3bot19gU75gIGNr1OaGV8VXJZcornIf9AULyKPCh1VDY
DabQFZ2cKx1+kiOq0X2IP2lz2zlPwV7N8CVwoghUEbu0iL6YxfmCNExnbVRb9YUn
TgRIFq0pVSEavSyu4rFa1QNFlcPghHDwyBxr0vNd6Ul4JhJjA3t/FHwEaMGAyU9+
SnZO1rXLSxBvajLzhOCzhYvl/2HfDd6cD8MCxLnZ0y16s/LqDDtFQoXraxdmyJUO
OEFaQHcp9vvO4ukWClfcjt3DMI9voAMvoD1jE69pitKcPXGlUPuvHfHMdv7Az2GV
33bg8UARpxzRWinbe+IX8EpPWNVBLURTyjPE95itO9PgBXWpUqD2F12Zx3SX+tkN
BBAPeUWtinF9zvj5HEUjt+hByUXDcVpo/w/mbGYFDbD7jK3pF1kAYh4OkHTuusnM
r4A/BeOMoRLVTs6xVPoqO+7XijAHRUeIPULTHThlIwmpda8Qy4RpWWGUeahmAfoY
IE+YI+HZAFINekRXSp8A+kbsmx0LRpXg36zFH71Z7/UQhigloAvyBydVYmWw91nZ
KOvT27nPI8KxuUCrHYB442OPg73kUk1mGMWinrxvWcIpjc+Pb5XWIBMKMHZCN53J
cT2ncKDdOeud4v1lCs3DeJzHem1AcPSZphqKog+wVjdStiOjxVLm1cV3uMKHWVrV
3R0juG24ia9tYhroKk+c9Jq6q2+qfoUzI1C1C1xo/RcClhryJn+00/9KUra7Cqar
KXb8dac6IkYDM3zBgXaKqcJtVY6rkiZNeLHHgSJyn3SfguxuX21YJNS8uB1a1UQO
8Takmt/9SKjavL5L5gROG/NdzuluWl1b+MWS7iUUhDRGddPunktPu6SAT1c5xWPI
T761AS0yBTBawiAlPzaQZ9wv+7B2u8Jy5XjZvpgDQSX/CRZpIx+4L03RBhDQOPyK
NkZIq3CAJH2gir/Xfu8c3nJkxxfP1ifwybBQeW9fHMKNbuFJt0VtHBkQaKumZOLh
5KbvtMqim601YzFMWoxp7KRogTEilevL1gCsQWkI8nQGWRshKgdap6wIPiD2H79M
TNESBkEdVUjnWHPVBJGJFh0JTG8YBNC3OKHURBJHz/YiYxuOqPsHsIYPIE/ZIG1h
`pragma protect end_protected
