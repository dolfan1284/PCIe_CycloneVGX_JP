// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:07 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sdTd1jXUmeBztoZcyhIQkXANvpY7Lz/SjSknWPhZ4BExjSjCH8raAABw5OCNiu++
uiwFmIQgqp3k3PQMvPN2kKw+zXKAqtKmhBTzQD/4MuDR7E4tGp3vS+EVxGaag6Tj
wsJq5EXl477NA2IbZ5D3/eynMN0747OQI+23NnypHRo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
MuVdXddUgBN896Txu0lbeHx4XDEFSz+PYXYk6AauzWJCOSxa2NLbNISdtgU/nzq9
8DPAnhibBdakbJWRWiyHvAPuWh8/rm1dcEv/ulyDveV67wM5PysDbXsl/s/RrSrh
pnISnXWoaGgvsA7v6E9ev8Bl6IKicVdcZciQGXyySYKRhcTeFlHzSNs0YsUI37ff
oJcPnseqijzP8sDVBWVlckUuh8Va0vyRv7DtqTXQbNUNOOZssIfTi5UIbO+uilwe
jtJcQ/XGOtvSu9WMONyvIv4kcOqarKgYwgD7Qatx0XkFbctMENnox2gsyEJ6neOi
oFx4cghtaujE9J+WnfU6T3ZNcjml5qVGiiopMHGlijS762aFie1QrR/e1w5YbOko
l3vRUZg5VzhB3WDstuZT5LYC6uSCfPMmKlyvo/tjLDJdTqUqLQxDELQBhsqSutXD
xhHyQ5t5ZGq1PxXF0YIVqL4ElI5lVOFRU4lYOuKnXZP2Pd8WKRDmBkQprH5Hc/Ou
q1lzVA6q8INtsVWAakW+kiiv/fOleZv/8gp/1k3exDJkG1sxhycYYJYCox8XaI+y
Ols6IKaTXKdkceoCzW1ftErveAPauRYs/Ge/SfnA/N7V9Fpc4c3z5f1KSkzZvoIr
u6UcuA9FBiKQtCl/9Z+TxYz70HEvUlb8HXekfPz2d/yvP/96joYZDGOnr8kGb4ew
oD7zUPakgwHkfV0dp5xZ6hQ6omZ5mQ4Io30kDRUp2WPZPmt9fsgmWkRjJ20AhI2q
TWpRFArMugehIXpQSnHQm1on2zOdlrTwYKnPRdW7g3SnPnTel43ZYZbUgR3bqM/R
0crFNBVwIr1jVuz/QJ0S67XUIcr5xAjjYDZ2n9RhXOwz2F6HTi+RjJVsrpzPt5v1
RESoulYgpVW6TP9komHgfUx3X1kv35KyHbRGLurh57A9Mn4W57ByX0DwQIunMIkf
lpukl8wgMlWAlfjox0fBkYDb/ozmpz5Q61895EVawH2+SnqpxYeJaVvPui2QoFNj
QS9Up6Jz/OeQveaQksOD0QR/hY6zO3KMnAU+4qOee39rYTya7NAveGBStgROLVJv
M6X2VjpteJHbwvdtclW+Udclr/sFfyTtAEmidZVY3MdrVD0YYwJbhcSxxYtuOzaa
oPmh5nfEG6smK1NF2uf7B6V4GxKTQq4Ff+sa0xqOTJqdTFLBYd5ZGtOj7wJJO/BH
GqDMWgdn7M8nxbwE+5uxyTVFR9T9g3EwzcKgaHr2Jh0B68ExMztibmFuK6qkWqmj
xUMVwbPE+KwMhBXUiqJEmkB3kQkH1xb1hXsXe1jNNLCH6hDEgqAzRSGw33Ymgl/8
q/xVPclCa+PPGHJtkS99vs0meRoYsXuEoM8aQdQstwJ+BnJf02Pt3Ezhw8ULgSdE
G3oDq4UG2ZAYYlU1GE4cGUnM0Ifte85S//GYb+oHGOR7NVNFUmIHoSnEnCkTK94n
eunP/sbJei6HkJLGoyiMgxYf7cTvJMcHLCc0D75OcKuMJehdY2aW38NsgckuW6AA
QTaomaVrk4+V6RH7GS3HK5NjTaDhu2R1jfWTsN28bfBj8y/7+UZqYY/7ACtVLClX
QlZz2VHh5Xpbb29/tS6lW8AsCXVydEUnuz6fCFaMinFjZ6kh0c+DMM1b7JuWb29/
6X5azdLEGzpKEmDFjFwr2C+c3NzSj40I3Sf+BJSANhr2uUc0JLzhg2gBwV034J4f
7qE0twqw+TRghlkLx5hUEEHCJI7szR5FlRW8E0g1cYTnQ2SNtVyX5l2FpxSjyHmX
lAjSoU4b0SO8FULuWXUixR9OV4FkfLO26ShyQCn7PUffoWfZ01b36GJwOg7YdoY2
z+QiaMMiiTg70P9wqeHG9FhQ6nk3MrVuJhCR28UoSh3+Rr4hmAWB5KsPSdE2Rmim
vK/ZiLIoSrw4B8QVL7iix36AIbv3dT5Sq+T1bwtXs0WTiM7ByLta7nmB98EpAaAE
FIrivcBMRznpbJaXlTSUjDwEvc34LM5SmgzkWJjCSq4z+BJBuhwW4GABDgQ7D6fn
qCqXEwybyY9lUBXzRdPpzxF6aeiVsgUd7KxZhBra+CXIJK9iwuEHc0nA+PAiTJhE
KF3KkRGVSY7eE+ANxDwu3ZSF+/lw8vncM0f4ZCyz2+47UEZgltqmJAKtFOe21dUP
KXOXdo3VUvHbj5T9OsA0ito7bal+jtrYiSa25cazEWcV/B+OFKzkJiAIclKcqlqV
2N+YPnxm2neOVgKr98JoJ5ZxvLsTQFb8tSsWeakb1xjS8sQ6tAfYmpJMYV/Cysj0
nzhSgbqJ9/2rtmchCsxO3Gn/hZ7va+L5B9rYKEWmy4lSLQosWDLwxSaO3yAUjd7x
DhL5xM+AO9Oyxpe5yl1bT82N4OJfO87+4DDBlsXq/xS8JbhSBoibSzBBiKNDLJBb
VDgc3Cc4INC3mxeF4FoRzXhEHKygkzTCuI1+3bIBXaXzR61UB78zqIcLSLCsAqBT
9KSuGFaad4EyMJ03/M7o1kdS4GFiqRTtnmujuK2dspPMr7yKLDslTn7mXxS1/fDR
zBDHg1vqkzJqmHYv4FfbhS0nZR54hbfyg649BHor/2eNcSNWaaxFsMW3oDeKOzhe
RaHZ3UQ15ctlN291VX1lqxEhXBOjefjtXCqzex4fpB34FHqFZz03E9Bu6RLyDs1L
KdByRjQtfJ/FUfud3UV6LgGdWv79rxQ3yLCaq7n1CLr0KyQJFw7EkHMFx6ia1uoc
FbYAcl9qK5Ke8+sgrq2eXxhieC6ov451hcuoXpxScReKqoVP4zv64zAblQVvVa5u
3inyTuldb1s2OzKnNp2xMSGLP9sgaiaEnX0nEMIcSY1GUF10bcvIC8iedwVyTBm5
t2uBag8X4RuLfyEQo7AQEhQdCAQmR0NY3N4TMCfPbIIQWziA3PLKA+R5vvoy0q2t
H9nMxEoAw1s6nPT3rzYU1IEHOmA5JbHZhP18Aa7E3nlp4/IkgY+qnh/1aD3wVB4t
8MYc91VQxVYANuaXL0OoC/dqjmL+w2WqMSEy7/4p5GrplmdFADMAgsNrxlBWV2vI
Inxg2AltIPXkIkuASNusJMqbzfM1g55a8x6JSEC///EsS2CB0r5av1g+wtCBU1Jh
2GCuOPBFoctvzNs8OzqRp04qFcrxBAAS1g/IsQL6tGXIGoHJMd6dAhuZH1V/6Gum
fmEqCs/LKEMNWmwZJun8LqdS/LaF4lpwsHhGe/Ky8FK5b0mLWHtU+s8lkIqSZvvF
zLHRlroJoYsUCwTaYKSoZWUgoyv9ITLZyp3etzCWs2+X/t21wsZzyV07wEnQtuFY
gBUZbv6QLeB93TNfAkpiv6xjsZ4uy39JfXPKOfQ2wJr6nOn3qu4Yrv/mKfjKcwmp
3UPbYUGJdjSp0sXB+nfZ0ItJ1E+qVzJcUa3T5KaJakIfNNcegKSk6HxFiKRx/Tz6
ZLPkuTlCs8spW0BCtal3OEBU76qQKcX6XflcbZskPk05BI3hSv/kUrG8bAvcHW5g
KnywApG43WHPbReSJ+hMq2jrPaDRL/JXLRcDtxTIWeAbJziSz/OIV50C7MnkhK1j
t2g+xDA4GRpwvVyNGHIkyEmwe4nUqlpdxn/0/uAm0751H7dHJ4ySA9NQDemRPHCG
tEvTcklMRosL+zSUQ+rdm7PEDgf7wyEtENoMoqO5TxEnqmlA1kDiiwf6tFsu22eT
pTSAcqR2wwzyMtO49o7hoT0H8JDacxEK0KQ45SHa5xHz4sFH6pB+Rh97Vuy04f7v
1oEfOODSO34p1XQTiESWOLyvXkC1eXO8XNg8EnBcWW0h+zu1wv1X3BvO2cTOZ9gz
2UlaL+pQLbul/OtcFGgV/za7w6Dv+sT4RAr0x5gdOmHltzSDgYGXFj5S7jTpLK0G
AjBEiOK+5vToWltdGj4CtW3iv7Hyb90MqabhytPl+maKsTWfpp7xDF/rfLTx0x9U
x3hUeBC3fJpR2aiIJu2zUv5fnA/q3iOmohBny4ANdgkCJRA3QbPgYh6yWiapvmbt
rtlGkRmJkJAlagTodhpWr1RRt1pUQwHShZX+R815qBDcNAJGSWc2DS4aWkCCZ3zy
p2p0rp9GMldGV/rUHOu/IQclfzPORjE9ervXOCpQ/UI3CwmvJgLmcTWdPz4DTk53
INV6EXKKqVQmPg9zBOCQbaqB6kgkL4oeDWj/ecOth6jHIcdN9Cwk45z/5FFsdt1U
2lKVF7nQqbcS1GG7Auld0SieZMsIMQkFNoylbbk+QR0K2G/htgr5m5XzOeGySV0L
3LNrp1XJqBYPvhtY6smpIfx16BArdeBkv13OxT8XM54/Loij+QRf67HRMLGx05BN
sXo9zqL30mEJ8mEwnpLJA+D0q1hAXqPLAVgwwV97ktvKrFP3MnW0MihCfCWOTAa0
g0IrO1J8L/xRz00vjbu4DYoCButbFc6knXt7wsdTQI2sfHD/5k7hvhwdJfk9OQYZ
02/AXO4pFpEozQU5OqQ7s74APupuQi0AGBVxEJ/9rDz3Gv6nX14UxNfJcEkmW5uY
uE0Ys6NaCO+v/T2GW2yKbSMGxJJZ7qqqlfOQW3/0DFnZLFFRO5DF3jkmEUbP1K7g
4o9N3fPm6TGsdI+wo/iYawQ/4jftbIXHRrLrK91JYTvqkP12Yzx88NbbPcTNYHUq
7+woKo14xm5pA2WE4S7nxBYpUXHGxR4f6PTVHeQhBaPNQP61YeNC/Z6nnYm6yyAO
qU5OuPWGl8+aXyVIRmqMzHIPseNA/fJ8Qoobc19IXmdy2Ye4RNSi02s06Bjx8llx
a2PUn/3FtdD8gSOiQxhC5WrkiavptbNqipxhgYuNyb2rPyr+ZBshED+0btp5wJER
bp17qujdDC7IDBdYcma9ZXYSYxIktr8SPAelkYKqwZorxM8W88DtKjHH6U/WJ+BN
fRnKqwuVFjtHcj+RRaIkdkqkX+a9R2NPm9/NFix4eLX60hbl62KjhrqjBt9+nkqt
1evFF2OhGJ3AkV11HhOy9x/+yxPGW65VvsM9sXZ2uoNqcHT/2SFh2brf9XoUVUGi
gPef9J+Z7peMdMsmOCnT3sZS/I5ebkxRy287Dn4kjqQ/cchawhnuVSsmIp1Or7Gx
dr4AeXYoWHp/Jmh3agd/ebcnH9Co1VkHZbCDjpTzKitpG4L1FWBJzo8med+BR6ox
dmn4nja+jtf6ABDJcphgB/CFkKmNNlwI+xDC8ODac3F5AgcgxdxjDQeiU0qbtdDU
xkt34Btn8V9H2dxdjoYYd2nJMEKPFcXemJQ9ImY9ni3XBsJFb4QUUbDE0NDiAcOy
/F1wT22KK3uuqzNAXK2747h+f33osQBI/4GW+zQTAJwYGbCNDs4nyMGrVxeTZqAq
8rJALdPwk1Eymg/P9ov6JEsaopHs3jRvZy9kwujZHc2pJCoFVWPHEOez+AGdSihz
WbGQ4gHfDymbFhExrCeaVnfYkuNN996LQ0F74FUvqQ7FMlgOEMcmsjiTFavyqTDw
PuY9jzkQl+wwBPA19sieIHt5UAW3uYX/dLbdYcwywlHWZURhaXssxx9xI+GweAsu
4YQr3KiKnxeuVgBUOhIzmy/u583K/FuGrptUG8J7Dzh3Px/dNtjQytMA7naOraw7
lAqimA639WsSOyshdSL5tVvygdeajZgqWjeNIsclRDjWDhNCVe7DJm4kDJjn6zG9
+1Xe8BneBZFkJp6CL4jiqX2yBE33c0qESkEuiqui2p4F98Wh8tUyamOsSq9hbeFa
gLSOlGP0kEj9jYnAHvGDo4eUoGg0uRuyn/a6VbK8b21z4t7thzHqNlpcBLc/3u/N
Lj5yjrGshsQGhiw/jALfqsShMF7KCXHM4HmHMe9VyIFhIANwmkZiUMoEcONwdpKK
kPyQRzP560HfwaX1zObchz+Nggd+MXXQ8hwELZy91mvW7qepZk2oY827EtPAmyy4
oEODFKDbSWjD6KI8baSZsj/3sCgl9fVpkYyZo094WD5AFD992MPwkKyiKwefNDVi
pPKcq7Y6rjeX6N9wQnn3Jo+tKFcNjAr1yb4whJg/wVc0nc5Y5GAbibz4MOSu8urq
0d+Fs9FB0fwKR8vOglRCbFxWLWaMK6Ogz620KrpbC5aBimLkH0LBBghHUgj6b8Sf
p81VRGgSNfbHWviPsPVk4dyOkRvwYQZothFMmlewK97MFp24pnZM2ljw5LFbTqiH
9IJKycwq5+k7vV0pinJZr6olvrksTesaUaDvZ9ekNqJoV0D64tYsiyR4Z4jslkBf
RnKRkYODrSQJJX7S7GcBMs8Z5cwN4LtU91sn3LJcU/Smne1Du4/6Y3RiSsRLgt0u
d6vLnauU40BusaNfXgpBqi/6G8IJwz9jmMWw7PARIN6OFsjOW946P6j79/D48XCa
0DfgnQ8DSu2KVikb2iE89f4jItiwOQYIQ4BxUFkPIUrq8q7CFcuvJenvbmLI95Yd
aVq5y30hiYvEUFUORgFH1aJiWvFP+TD+K45Od9wu2UzCCSyEFYe+L7W1rReuLfSx
raa5pNS7F9bn7gR8Z9ryDagDa41a9d2gv/fT58O5t6znsjPaEKfvD4SoeFNEwNZL
U5CAwXOX4PG34UegVEZiI4GlJaw+klIMI5OgkAHmKymZdEx9JbPF3sDFMj3pmSzc
NCFVHO1bAWDyz5qtyeiMp+sAT8v6U1dyzdSX2hJv1bPOvfP9XwDkd6F2mT/DpxJ7
/nVbzurRp0djBCwTljMTc1mIgkQAC6WV7Hx7F1rkt2/mBbmVOxNptCFGKRzHIeC5
Z0dyI9IZtoblxanICVELeYIV0+gRSMRJ+u5nrbBrrnUvu9Hj9h0dLbTpgl48Eftx
0/2MB976d40GF1h3MbV7nSl8ssOSYLrB2vVNbjhvR7N/6LDZr3Mj2G/ESnCD/BsQ
VJBiyCiGLgfQSmm+XraqjnHLxH/QA+CaM1c1yBL8XOmkf/nnE3TYQVcl5v3co3Hr
LiZgKixatiOafaTYtQ053AUEeAbX6+IJMVMj0NNH1AjHU7sDcgRhH2gI88YMjJav
5fGsHbdVqw/w+OJsqbXSOmScB8aR4q4sHaILbClcBaPsAfjWfxeuX1ljbjP8WRru
3vizquE4YItk7La/dxByPhUW+CqGDg7j86RYT75mME9v36rLZ8sfA74Lk3YRaSVr
G1nf40TCn1vD11LiRWJXeeWGZXnL0ptjXaiURKABlMDAoyM/uHNO9731wImeuha4
LV7OXWg0rPmAbhBFvBuasr5pv2zopFqNtJ1OdytNYL1XqB9JCuWRUxKCJ541O6SB
F+gvYl5v6DCimo9zUamYplKZdB6kk7ls1lIq0UGWhlqokzmmcIPvU+KiZ/bsVMZG
1RF55Wr3Ic9Ne4cWfc3JUPKT6LODFG6kB88nj75CaL0RyZtnPm2ZHgO4WmMfqaie
w0/fj++gSrw8OFYV4Xydz5eD2QHx2TtFJxkGMS28VdveHE+NbfaqiTDfqQuM9jjw
Yvu+BZm/7RQQ+PS1tjFztx8+fAN5QBnDSahqNyiGZPXpUlK9bR22rm0mOiZgqf2H
pGvA4fsmn60SUI6w6klya+JBPD7HgtqAgRNev9KpgN35WEzY8gPXSsa/s9m725zA
U3zZTJd4gAiq0f6JxKwyFMjYUsNEapCuwlhuFz1vH/Z7FwnFjXKn4K2o/Ss+DxX6
J3OIITWy7U0DGUQY3tv7eThbPqTbBZKhb/SEStTkWc5zGoIOPwwSTcBCpQv4cEPD
lTA3UE1Uh1+fB8Bu/9ET39DK0la9J+R6kaZUVEZVa+o68N84Md9SbQRvE1dpj8M6
4rs1IYu54Sbx9vmbLFX61JmzQrhurms/js7Y7MiGBrD8iCxiQ2VL2BUZUm3+UlOx
emiXUio5bWg7P6i2sGvxZTI5kjUMpCt8c2qmd3X7994hBW1s2kzQUuFNQ1NUSVIk
f1XG+BySeDW/Yzv4Kxg/sz0S40HorT9XOYijnQxI0KRSaxsbgOSu2GNKm/N4Ep/x
KXpiHskossybr9VXrEjJPRve+avGi10NYlUW7AoXnV3clbWGs76Ud5RXuw9WKuel
Q7u8P5/3/xr0VqVGXmgGwjWmpM+xlKXqzlL4RZXGsLj8ek3hjZlsjtfvHo2NIFOn
vYIiA18knGcA5gDR1lJqvtE4t378UFtTj+LQhyYxrJx223NP6xAzrAgOVDd7cNx+
hY86I1jEUEeILiD2Rs/HPI3PLSVJxUxPHc0T1IkR9q06QfGWxcVeI4Z95v5pDigP
g71kXtsLWfoaRrtxxEpZuw0D1883+JDB2PDiOMufJHYTkUIR6lLzkm+AF/exUN0w
viQzy2iUrsUXosgLF1FQeqAj7AgTH9canCYp7pjV9E2CP/RIkaxtk88AvrCsYB8u
Fff0lrkvV1LkY3wTFXffautjBKoEobV0pbRcpCnJkYe2J6EdJD0v2gYLntKWPin7
nT8fwDdJSNke8bRL/UWjTR9hSx8gtk5USzrDoIfP0OJilta8H2rhvWUSPlEsrg9K
wsUBekhx2YwgRpeCitWh41b9aLqdPMDdjVjN54DQ/c+x1o5VpvM2yhaJjf/mNu+Z
O1qXh2CxNKFS5yeAm08DTRsXkO7idHcqFk1f+JRKWLyPHP/zF3Vp/XaF4WeKbM7G
FJeI6XNPX4THQ2HDn2a/YFWPzAbVaDmZeJTHURPkN8J8qYBuZYgbBtDMhaXH2BIi
U2a/hSTr+ymEOn9eMaHpR5/XIhKtYVDnHw/9vKUzoV40UEvZQIE0Ko8jiHJxe7Nc
wqdwlK/IA1zvNXPf/ggJjD2nJBDe3ZGTcgwvo7R1EKHkY4EjLHFKftmBvm5UkAtR
CKL6l4OMhNdojIUqswjTYRDIXQOZHVeBW31KRIIcW0rv6ZMmOV76k38FQdaipT7/
Ne2B56BgKcwX8YR2HhOLISR3ZuZavZ3ltDG19cGZmB4DBnpVzbEmlsklzqcWTT2w
0PxOFNTnwLi1tInWGyT/Y6XftLz02dAhZGWju5nqOksPqeWsWRT4x9a+oH4Y3kxS
Cg7z3J8QKZF+wwwr0iVUcPCeTV6ja4b3M8X3xHFIR7+85OfYjvnEDa81azh7YDvD
7g2m3xUtbWNh0NuShPFA6kQL6X5BR9hyqlie/Yh8KfS4LwB/oXVHQ1VDFUyS7ccr
1FZNSZG/QJ75H8iWljU0/75uuYt9rmjIoV54K8W/cq9zQ/p/8OQlct5zIcsstqNl
T08VZHheN1mQPvSQSFcrqjDqF6WKjvRBnl5Ux9exa1i2YJipinkLA9g92Hc/Vywa
M+EvCR/5EkczcEPUCkJ4LBKDXkNB6U7Z7KdZF889SBNIdIbCWKhJg7KpapRuPSDO
NRXrMThLMjVTbhPZn+Q8gaIHJyORONT1u9zq3TDMcxBLzD3QsBx/MJAUIOqBCI3N
4ccJuNPp2HP5BSwTT4OoLpqUfBevNshGX2wdlNrEjUsId4vKnlL7p6jdZBdcrfh2
76reJfE+Ft/OdaXNcocpOBdTAITbVyDLR9oFJJli4nyqJbNFmK4x8HXMQQ4dA5sM
sX0StXGsiiPqJFTxST6Pl/Zw1lgeWL5n+7D/uqS31JFgZGaeTAC1Jn+QBI6lzFHW
UB6Kds6F6j7gmAGBjA9o9fLBzQlfGiZ0qP0LzZO0z+xfzNFVquSSwxaU6RyHyG9b
dj4e3x4n8E2CF7KKXafpZjJE+3gbSJ+q1rr+Syhq/ZxdIFVDQx65FGy0L+sFieDT
ybUZP14q9e9zKc76uIDUqRa/UKtTX1STwqlCe2X8xxReFq6gYSGUiwgIQlrslEjA
Lrm11k5R7Sm3pXqaQZ8lVFuzW7q09PByBJkMKYvP5PNNIEyIekgOz+34QfpTQ32S
OY7fYDqlLE4nq+6y5JEtluB9n/PPc3Zi4m5SXFPFb3qDsau/Y7lk3B02OREW49JQ
bthVMgieO171P9wlVqYN9pwgJ6F5TIfaZBGeGZRta+27Ywg2EbMZvDlAzTrmwSYL
9l8sKoYZrToScj8CRzTMkemLZKqidHmO3CqxrFWCEftR/obN5/zedQa9nHUC6+qp
pXuaVoOsyqct1ss0/zlOo6bwNIKw1mN0w64MtqR75pH8R0SRy4D6f5N/Vawh38hg
BrJBiyu4tsb5B/a6Z0gw0HAhYgIgSCYzOjJQmMuv5GIokvZrUh1M8ptYgbIpiRdt
e2Esv7OOTwaxQr6Pnqm8kVaoumuZHfhrNCjJoxHRXiRZjpCOJrA9ARjHGXWs44N8
3liklx/sG2z2dhMP0S4B7JK6kedYDohCDWIashyY5wGJEtvU7PC7/o1F8POkeprQ
r94dq7jFwBUxZstaD/AhCq2+v3b1y/05NuUpn3sxWY9HPZ7iHWm4aSOtjhUY0Ctw
tyqO7hKGwAvqe3uJpErc31tO+HsiGHigWVYf8KuOZf7k1BP6i2EnCwaNXVOpM8b0
YgJlb3TVw3qf8mwJ0DNwhFZrasBrYpc2cIJ1Sw4eqhj5COK3nxQkjphxMnQ/GZc2
TBy53sI7jyHJh9urmNDFltTKIQMCRquNhlv37tmX7eFrMtyha2LSIOWfI0BaY96O
`pragma protect end_protected
