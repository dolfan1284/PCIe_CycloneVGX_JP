// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:58 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hn7pLNVmwbGfF5G2qcq5/tIxjllSGdl8HAblpFL5KH0svDaxe9dYGS3J36rdo6lg
+1lNBc6hiSoQfakM1b13dB+eKmjvp715jkP7bRNpskQ48S2CVhF1cJwJUkb3GZdE
D9QV1w1LjETtANq58NKOuNsoqlaOcsev+BDU3CtU4SI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
daM/UygQ2CZo/xBJSeo8rJR4d+5hDF1bfTydVYwaupeB/S40seij0266boTkBmkv
6X6M8ozzxC+IZh5W5l63oqGzRSubNdMfD74xf0HuB4pTZVsMkrwipPVrEcYyYAOy
7dTS6kK58Ij+CrHvANkJcVkfmrRaxPWGoa9fltCFQWkHXG3tbeJL6QxZrcQ0+/7q
DeVIA7eXiFJenjdS5Ecz3d6yGWm+vvgIxfrNW8aRLy2r0IU3X9euA90qlfHppCj5
yRxR/7P2labdgbqYxQRaw0sU53+G/7SQJ5xcAjPqAZkEb6h+Ga9ANJOgGe6urigc
scwVSOmjkK1+GFbMfnUoBCR08Ucd+/KIKFr2i7XCLoQeOyoPEv071q5FLChBkboZ
U6uFQj5gXiq7kl7it28HmX6MIPvVrq/SQQisGmV/Yx2L1sDiUoBsxVmcLmbYiBtW
+DXEa1kleitI2pbzdeSUw/bi8Y8MNUrTUbOXVRg42Xc7tj25ZaLaHFNw8RpKwIc5
YiJGdow7i0m2mPA0Nwn1xFZpjHxy5O3UCoTtDRrR4wCMe1IPDFekkrOmmPwPvS3w
CXD+0QZeEvWpwmBZbQy2xjAEHJ8FBhHRsxvmvhxY41dFzQvcAf8D8Ss2thSe7MjT
b+TkFHg6howDplKQPwGYfeydYSdQYrH44e38NaqABRbXkbdexZ+5rWoRIrftqAo6
xHEqRKYZ3goqAbdWnWiy5m9QZ9QQtSjBF0lutjhKLYTN6oXPMjay2MCZbOxK64Zd
m4x3KTM2+rdlThA9IFltP/qgcU5dtHKxFZHMlThmvFyDPl7eNOGa/uUjHLdKpqFc
D39rq2cb9zRAX9x4cHOqznr5YOunSP3KS3eQ9J3tZW7m46GMnsWwZTIcUO/GycaB
aM6QM/10/lx5XaZr93C5zOveLYyUvwkHiNVc0qepIxcPwaPu4fA3PS55Tw5tN221
cpmAwvtxR6U7CpI+E5L9piu4C2bMGfbXwaIio2eQ6xGT2aYuP67t3YlN/T6pn1Ip
FDEU8upYdTj9jOsvvvGr3T2jGcyGGYVZLDOOxC6x1mttWtMr9wfKOSGRHu84JsCL
RQgX7HPB9JcT7FCzJ1c0fdMNm52Ue6BhmNCRFA7b2+2jVgUM4rYANfZHbvRfhj5K
TNy7zLNkgGqr69nOIrQlbNJ47xS6Eh711ZWSO3XXsB9UtZRuwZCro1ByHc6LHdan
tcZhxERbQleBHJn2oLK73NoXgvJfXbhKKGkNO+oniFk0wM101iMUQLxS8BvgI5zJ
rgtSbgbHxFo9eqhb0okFnIFafChnDJ+jntDX6Bv1K6SXstzN7TMiYTEpme7VhZXI
w5QxCKJxX4F9pmFRRg0Q+AMRG+/ZR4J57FzTAu+B3gXuC0taN9RZ2LgcKEn9DSUW
6NYp+2I2DpTwipW3E2N0yXd8RSjSRUez6LWN08F0jEFDR5/9+Cdxukm2GY9Adu7F
bU7Qu0JKGYF/fLpPGKnqA+BOH/dVw+q8L5+3fYPqpAtmq+SFKacgbTAduTd6LF5c
EYf6/qXk15rvUSRaiS8lD+oOPAQFm2C5EcoMvtO2hbL8n9fQ93aCyXDP3aUfquiz
1yKtMINBmRh6siRxPHrrOfM8zc+6tWBLBi6QruyF55WUYmv3XOpDwcybethRwR0d
LDjf+PWo47t2UI1dt438wRL2bQior9Yjq/vhF1Qu+QnLzQuYwdpOh5kDYJaNBI/n
mM50AKlZaEI91Uo+FE/FxC8njADmw6zBv5tHkjPrdaBAOJUPVP2hjZhi2FYh+G+G
byDDGCwz/LBZdHqMoHs1gsPEzJ7PPhZE6dgyTifXzfK663XMDPC62txZNNd7vjmY
cuGqTCNlOYAQJGIiNSe9kbbvxKfC9Fox+HXZF8eD08ziSGyzbr+U4XZ/NJbpcYLa
lIYYnpcnIuPnWU/69HK/tYJcQjBGEKcsWq5xcZqylQcYDS69speWZvX/sYSvR0I+
PN4y5jxIi8ajUl+jnQsm87gZjibsIPyI+ZrkFiRmDD/dJNfdD9ZKl+6C0d2Sctiz
ffqXiMl11E6Tqkix4xidjIZpSrLwPLmhrnJTVptDEqxFu3sMY8ZR6VaCZd9DbwFb
pkP1SSzl3NcEIY8XfedT8R7J7vxDYX9xEoMLWlPT1kmC1MW0i4CoJrDtH/fzdvYB
PvEMALaOo9l88EqRfsjjz8Qw+qnhPmGaECxod/ey8Dr5vt+LsL8+V65FYfPM58o5
6tTupPlczuxAqX3MF2/XYBeCeXGLPMW5pDayxIQJIZGdy1YdsJIVRamOE4Neqcl9
6M5rjknJheCahq4/rAFJ92RkvNpKL961r3FR/ztu9n/jM+BNb0Knfc8ezueab7RY
iXE599i+HdeqEGvg8Lkid5pdUz8Zul3GlZqK6hPMK3xwM+y6nA0DaOApO1rDKWq6
CngEhz/mh3iMFGCVQjnMjIgXm2JV1r3yTwS2ijGfYn0B8SS+8TGIbGQ3jOO1uB9w
gjK1m1gJ+Ce4uyIrnudAc1VlhsI9cvNy6iCdEvzlEGCLkP5FANLEPL+CT6MF9c9g
owsOIbSV2GNNTzxt8ZBVGm7ZO55xdtN9rBykrWV3MBzFSp99pvkOFhjKEolCVxn8
xlKAsoab2Xi1mmw7EiHyee0bcz4kUyeyninC47BdPZdmOCOxeDD8ApEx073L3Awc
tAXeyQL3dLD4Rulm3BeNpb4D7CJ+VG+o6MielOI7RRLOOO94sYJWWz+VHThwcebC
8RqyJ8UFkPcJl9YKJwfnfdTFqJ02LLLZOqJ1mrQiU33BGsPloobZ4LWBKV9WyRS0
XE1qiCDo4tFhh6g2Zq7PDJbNp2Yo/dVC90y9ZvvPyrmoUND/9WwmEi4hzcPHW/r4
sWxJT7YNYfCRZ1DVurSKVVg51TU3nRDCxLFqjTAZiR9wmoifO/nTrT06g7p/8PzE
Io1PhhpATbvowOcxLwEwBUvK2VvoGBKoJKc9HPLDCez16smFw9+geLfnhscl8jl7
KXCuHP3w8gI4LXzDzHri3CpqJ6ahswrg/FE3B/reToorvaNntyrkGppWwbukybAD
Kzmy1C2QqbCWisO6Kauc9/GMPAbU/vDr/NzxK8MaAO6LLoAi8QmjdzakLvLt0ePl
DyQ9orYUQ7UMhbWDYxtzelg9TKe/Es6mTP3PJJptUiQsc19wI8lZjqzx0S+ZFIR9
5SLoRNDnlDvtz9/nlpfxIPEFIVxnpCPPfpE3/NqYaiDgedMLa5mswRsaeu73xQpX
B6mlVkSDrRoiTznkiW0YqSvjXt207x2xo5i+s/APi73Ts6ZnfDbdNkFaLRx5AAYm
iFTh1KDrJr1aTdVCShr3ek+petE0F75tU4tJPBMuGlXWabicyYQQLFmcQA5+Io3C
ZhipmxLjonhraPD3BKi0aU/0B4WONH1XrsfrxpgDJ8eKdf6O/9NGPcbp+A2ChnG+
S95KP4UgwF+W3JDXJ4znf9LoicQ8KBbPbWdLy7RAzk4Zfqm979ygn2cV2Awiy5EK
DzzG9ud7os0DFjM77vfAN9upFpgmO8KOnK2kYB+naX8FzA9jXh7VIwF7F4FV/oZF
kFIRIBPnx5nfHlNlYliT4EdOS3O4azzi4J0CEQG6m75NSlbzeKwmi0oBMAs9fPr6
IXrvHP3xwkLgd+JeuYeiG6cQuwyiES5XeOFh02cyW1aetG2jzauFL2Yq8eRNR5eb
En9DGP88QIxmpEu4TPZgxudSBH6RMD7gZKIkTpDxyTYNK5XIrG2QMZUsSzsaYPhx
V5dMiQjIZXhDcuExk+d7c+n3zXwV6dfGHhPhHlwufZtRcxJPDuhgt7TtaUnJKPmt
6Sufi8WsLHdMQkuyRocYjUhkZLk938iA9YyDXjWv9/LlfKAm34L3yjSQrC/k0XHo
GIbM3xOYILc9YnZOiwVrEHKAgYvftDesjbTSN+I88N+56ROnjoI/lijrAQnITFXa
5/mQ7XP1XiadYNj78uMy5xObzMlqxNWa0AJ8Ya6Pwyh+RiKPe5RxajIgiz01WfBf
9cCWt7xaQ643UM4jbsiupj9oIvl7YPjtZpWxGMRdylc9E7/PccDIXk7J5sYmruuN
0Xnlt4b/a+XY2J2RLdrw4mNallf/ZbsBm4oXjQA+TVO/uQo7iavhUryj9u3U0YoN
ROCMWdnes186k8lKsuIaKz9rol4Q+V/yBwr0AFw/fO2N4ht0qDDcLjMrtdYTF1e8
sfmJlHWxOX84W+5Ms75nfKDGsH9khp79MiQ2A9CQONeSioNa1c8Y/q2ouIFucN/Z
8YdebNsrxlZ/sWSW1iFTkFahMhWyUVFr+YCwf8YSGU4hijey3hotNaRAROp5qMO1
S5JPju4kIh4566J+I5nX15f4wQJs1QIn+VT2YTrHkT4GC6liZf1hbHMtr5zlMClP
6vQAHApu5nyylKHNzn8lThWIeuXaIuZWug+pQu0xv45YDc/ESkhxdcfDDNzWWSUS
Pq/h2/jWK6Dhpkg5Z7r9A3hIBcYPNFaau6V5SOcAmHNA+cLajIMtc+sRUaAwGdYe
FtlwfJR3BQjfxGd5ZN+7zBjSOsqgEzngpZ5WpWIEHxzs3heoWrj9OiBYzS1xGEWm
oWekpEQ2vUex0hZHCLel3vWlb5Azz6LTFc68omaCO0DOt8KNXCF/9IoOtt0jwzz/
APOa5tL4kG+1kXgRNXcpwgqV290PoZcqO8oNbIwu8kmQJ0zIoX7NpHekjfBD9A4w
9f9dSPSkWU52Tg7pzB91l+bAP9wLuNmd+T3KTi23lQIZ2hkHNAElvAwDCoweoVOa
a5QseB4UUv5orhKVfu+jikCZx2xv5gh8Wz6YfiJxrpmtfDy4FMSI73YUdSohtlNX
Yuyt1me7z4LEAKKBYTtxKTa+zPc1F9S3oqMd6pc57rcBKaj9B3VonqfJX4QiV2Yf
TUcMhqS4uTth83sEjbzATtfprrj6LEA6oMyxFARuauZdFxjL2PiZZ0EFSiY2SZpM
Al82LgWwPP680UwYu7uFufjDbmCB6FV6KgiiPTjoo92MdTwox9iYwkpYLxRWAQmg
Hhp4EDTldRLZOwG6WHFlfXV07i+oMkSJgGbHIHH9/2Yg1s4ce5bAoLXhfsvfAnkK
6tRKg8bWZiQKoaScdx8RUBxoo0C0ybtJF0OillXj9gJDkOc5lfzcNEirlcvAD6Kc
jlI1oRoyzj7IqVVePFFbiBnXkmsmfRGIjXIQY4ePE8mtHlEKhtcnXKP9SXNdtXKk
8nGkYFKo3rsKC6RwpBOjMxiFlcIh6iJe69CIndsEedsaUY4RvP7EAY0O5AIz2zXV
O3EpZhhpa0thI7SBDaVe/s7xJI+KOyvb6No+SO7vVzJsNtdTTVGiXOxcepYDbHGl
lyB2+T9CCATmjDUjeg8lBKkiwlQoHUmAHdefdn2Mj66mC5OqRU1XrAyOzRrEqu+q
TM4NRZJIvytYc1qD/aK71RRIId/1joWODKt2S5jYv7vNd9eXvQDbwOSvRvLj2Re5
S6p4xCYUCf37M2h0Y9DPSbbr081ktnNPT9ma1EO8kl9nmOazPm2Ne0N72fzMcRaR
kMccYRpYtzaQXhE1QvNGUDPVgDQUkaY3rEHq+W6fRuSHeP9glBdkalio/EIdcSe1
InsBlgtIdCcV9wWlcQfMNXcOkKN/aC2akzfgVzy0qigf4znozm7fbLsiPAi0NS6P
2QtfHJBpPJPv8Z6kRFMjG0Z2RPUvfktuT9mHjmWpaQlWDoLl/tU0AFm1ZTJSypAk
s4Z68nTF5KYM41FomYFNJUhSaTbtg55z2kvYBj94rX2o1sNUqfsbbWmq6qcvqzMj
4Q8Ngs7u0B+erkye1i6x0rNcBu440f/v8ncTdi+tZ+VLDf4gQe84Sf4vo93INzuR
AoLc7r3BtS3oF1IIBVaT3eWpmlasatXmqyAlCK+wh6JfGuJEjYfInwvUtBPZiiOM
Q+yDv77DW8UsDQEoIOHOiUKNLyJRy+wOFJ4AFGuLoT/DajSoOQJq8HQcxQuAlPrg
ywpwfspevHr/GXph+SnG6KgsH3cmsWSzmxsMJrW0Icc1r6GjwRey+0SozX13hjOC
HI2W4rVpkuI71QVY3bFM9+6Ch0Hx/qCXs4pegcdFLQjaU36YrMXCfgkZcZjQ/Qub
PmNjXZLXzC6GEnXphl/Dbc06MmVQhrcICyd8DoAnn8PZuY1u33nXGodIzXUg6twA
xy80dq7qq8jnTMU7MZ9GzWOHj86AF7b3xOVyF9XJQZ8W06XiLt0xLpkLK8uS3y39
LB3A0BHZHkeyDBvJV51Aq+fHkjW2vb9NeOuy0TEvc0tjEGG7C5q2E1fBk2DLwN6k
WuPTMV3npsbluE+VnJl2hz2vVZi8UPOWyS0+2RFS2jv+b7sOLckrlgNMsAsDAm5c
GJtSTt1flSpL72i62I6stpqMvtirvQCPeUJSKKXCOBuB00u6xDP34uQYTEZ8hi0A
wx241Lu4aUSaiVqVVIY0ONBT6e7SKH+LoaARduEm5acCFnpkceT5Fd/iP3RNh2yG
+sPEr/DF8LR0uM85uLVJq9MtftfkaWE/g5T4CUR61/xm+tv1AhMd8PlMN+u0DBsP
9AA66mu5J4ZOmoEKj7+UtfIJ2PLZonepRVMI4Y5ADKCDxIPTpkYj7qsgSLKkbtA0
ItkwhDJfPYYYNTTHGRaTy/xPSiyqzN0mcI4Vj9oCMJo4Khf3YNmVjFfkjpHLk3me
eG6K5jHsbIj2eBNI7rwUp+p+7s6c75/fvuu8pw3amwMTyLurM+gweW96yVFOoXV8
l40iZuHHTSX2/WBcLPr6fNAk9vLo2DsO3oNKmJZVLkHzrVwAy4pf0njgiaTanTa9
9D8u1R11gkTmtFFXuOFzfnF0fy8+inBrrc5SvwT9jjofPbgpaZ7VbNkqvvLZ3F/i
NhHpTFPJQK/fEjUjs2YGhHR1uWAZEQn3u2mLq/wKRoesUpeu5VFCfgRAONmv6FZY
Zp1HxeXvbFAIVvLw/48PSUKU37Hd46I58AaT/tzVigKIFSaOyrK67q+/gT5qrSJk
MWGp1vwgwolR2fLr1uarigKTb4R7Qv/X8D8lzkLydWKtueH05HLnvi85T8uH4dTy
XE9sopBNAZjXXZ9/IgyG9aHei5J8Tf9MHIkK/hrieSBUuK3P7aGdMArT9NbY7j8N
4SlK2KxqIa13A/ApvORUCebX/A4TNEICqOlwvsUWS1/5AMeXS9eMS+0HjdUh6L7j
O2eWEPewANl5VNESTlQXx2l2Zty/MdGDFmOn1XzHMUkvsn878oBkHbC3cgE1OQnU
U7FcguHBJWwpKf2sXTIW5rTOY43IRs2VhDd0DQMeC2YSZmzQzvv7fKDN5N+VD6bB
7QSP3nULqYvqrkcxWo2GtgG4nu2mpInmhwdQjLou/D9pOV8zj29KbbaN0wPXsofj
FLUa5oX5pfgt81pmChqOMfCCxUmc4G5Fo+R2Lv8cPqzrT9cHh+zuIPgFi4wqUbIu
k+UMM+kUaPyb5jvxQh7WeUXVN+Z4rmQM4gkJvS7xDH5QOEVHO1YtTVtA1Rq1Lfhg
dFINXeqow3lFntIvYA5GYPM/iRJ8EdcXAT1TkHpJYwurn/LlpCbwuHnp2Iwb/fzh
eK6rTOd3gFKU3uHfaeKUNVGUKBa+X0r+bYCFOD6Jwt+JmBpBU0JNSiCqpo6LF8+7
LumAnRqgrvMnT9zAfmHO0Rx1TbdH51wrvmtE0pTQQyMWM8yRSOtLQqbAc7chXIC0
vcOyk2DVwum7COBX5+X8DWHzWpptMI6oMGg7aSBfaxOxMn5JTGnBqbMBmNI3gXXy
0cR1bf7CpKXlCy5bMqdtPjbMHzQrsotfbwtNFEBDiFVW6Hrnl9elVR2/i5BDktlq
I37CERsfetvekh7nUSpvUX5E9cZS/oSgHib4M8aSvY6sedRsrMLneqFM1oo93m6H
Q8OnJARnweG2LSnyX+SaBb4HdQhbpQD8ICnE67/caqKopDzWS4RLifXaTMTVpHXY
hbFpCczUWtN9vRIEXO9hXfsXfjmT9ypOzQCsxf9JMGw/HC9ogBWTUWF5y9NKfT90
LOo/wbJoAGD2JgeuqoNl6m67GxsmtEwJ2tLoihlvgkTBhLmdwxOzZstHPMyveAzc
fJSSBKumjLmChS1MEHfXi7nyFju/uCaLesC4i7jGHf9xs6g0nBbNUEjy7fbcE59I
dNIehGUxYvkNWm5BhyZ0/wQFb2ZfRZBo9WEDWcuCDcWIAyD4jSru1SWXB3WhEFmE
H/tjiUtecmO2UpT274PSrnUXbFOYB2iIR1p+Ue4tGTSNUOklNJAadwr5/rMMbtD+
fpwy7iwLadbXh5Q5jFfvAEYHg3v0p+Itg3/9N1k0DQLI2H/dkzW3ly93rUXx5u6l
6GsUfAL5i5f+jdympL3PjE/u37OqCs3jwrtC64zcwGXZFXpPSVIipIF28k6Hgo4O
IrXMXbDkPL/vW3EyXqx8tv1RmtLF+gO3kv/WQKUM4NxJLsxfNMANcB9N3etDbbAe
Yhf6ubUrS9aLKAEh1CMNu/ip4Z4xrIo+EHpA34gF54g0g3euZ+0BIaV4VEID4ynE
GwmyM2y0327IF3JECEExwwrGLjWe17ZwLzK5kyfriysbe40aE3y4Vtrb/I9xA4lh
y8OBulanTYH7sa+lOQPRcKIxt3rb5w0gf00HaBiZah5horumvt7vPhqKJIKzgYad
xOe73oBqOmM2evyxX9M8Zl5QFYdMvdA8Wfl+h0HstdsQoOdpmi54XQkTACj2LWeh
0aCMr/cbLL1reR2yzB7pc71vskpV+xklExCWE2cA0wx2OJWFmWDnLY0Q38z5DCYz
uiVjpgDomc1Pw14S435O9yYUb0NLNS2F6aBWwymj/uJ35LDLB19e49114SClDGTt
dARh+Or8YsKHK7h9VLaHklPheMEODBhqA9kThrHt2mk+a3TyVqSyuuogffwVJiwI
fKPApvFnrNndfzqGwKf0ieLRpOomwlyRoArK63yDo2WvL5w/dYNyIKS+Iu8jodaN
6YF02xaa/dtk6sDiXC47ia0umKW3BBUu+5jA7RN//mLggBdrCEU5exrI4NZUDdXz
KzbBf4pW1lLm8hRbT9eK1IwN7QchOwQQswAvlIIkrihZZGdqx+mYJRr5Tybf8CRt
V0JCRuqTjqPwn/4p2l56Lj2Y0yOZh3+AbbABVsF+Wx1VABHn4lsfqR+RS5WVwnh2
7UGg0D51m0qbnW40Y2XzZzejIkatGtxHfeNGcJylsC6RmuQVtvoj9M4VZyCLBqk2
ta1+6gJ5pq+32FInsPG+hcu05jB3G8y+DIhm+QdP65fIIvutQhohciKow2GnVLXp
fBBQH4DiqZxapM4RXcpkkvxhrFM3WVhN1DOBD3NyulAjWWKDJMZesLSKdA0pPwVz
TuHjkI45QF80H4fiCKdJR0IbplNqW2OTkbyIa12gWWeruYH3H4kIVK1yIprOrJzY
pAMgmqWVqP1grBU0GT0rOkCQ1yLHmJzD/v7d9nwOf5eiB02gGJtwCXhN4vmLhF0U
ehIpQtOvvmAwIs7pGquYopO+hlBUxv975F0LSEMYvDnQZC64T8zI/CBHieOf4Wqn
IVsXWIpQCMiR5mddA+8Cz6pzvgowK0SZ4y93cZY/Tdxd/nMrSs6wroTSiNdpXb1o
Z448MhloJ1z5/HMyVCh2ecz2otsZmjccXElFC7epL2czB9nvzXtX8epIcKY1+vW2
uT4eKc9KmgFN9e7N7zXzENqn9xqU6yK2EeYUC5Zs0uU/Q4O2aEp3QusdnaMLsKc9
RM5N0C1eaoohFbYHZ8t69j7bMNILCkbkzE20M2LF23+shBxP8yVsydgaxaK+gvWN
upJ0nfO/RsyyHTID7VauY4lesVVyg282aSCwuEhk6twdA/HPkbZT+Sw1LmII9RF0
2Hdbktoui1wkpWiupWiU8v3z1ZBrEcaIrT2osFgn3djFBMQkB439s4d+vcEjQIDr
Z2P1+WjCOqzWND7PJ3MrAjtS4JnWr3x7cJFeNk2+VuuJGFSRb7S1xkY0LDDdKyJG
ZHC+YalGLzjPZknRNkP6IRB+itlL/M3/5WErTxg+hGHV9GmBWdlUFkG8rFWHqMpw
FSj2OH+/8+dKBAIPdxA7aoZHawN2Q/S810n/sXGbNpBWLywBEZMC9WH8E2QTn4GR
CRYfaWYC4+Yubzanlr7KejycDjObYehw6qlahQN6/IvjRzjs4Qz8rHcL+Zw7rpcM
ykG3yVyAUZcy979ag6rFePfLkVkCchTzloCMsYUd9D+8uTbzQi+22UzFPKdh6bdZ
mE8E3QfejuY9ZSk3QgGvpXQOByESS12LCZmWGK18gOl6PdZEbzBxku4hTZn1r6au
R1HiQOTD6PED+vDOYjR5xKbeuNee2BSTmyvcX5nysu9YFfltywFMDtukHhKwXiyQ
d2cBpgpvrD24lZrcS2Mi2lC09oAh862oxK1hIW6cf2Z4rN2/ZT2FKGf6jlT8cvk+
K0dSTg5blcWob0CVqYQdYnxlLyuOtkHzbov2mrmqcvav98ocOvjtfdIt/UbhTren
Rk9HbpwutHtIFuOfg6dbjd1UxpCC4V5Gh8DYdASz1d5IYxvssLJB30Mt8MM9fwoL
AVOgi+m9Rrd8uoNSAm0NsN3xtljEOcdikU0sLh/xE7Nwx9hyMUCzdc/9jd/FST/E
fE5hsuhqI+bQBVHFiGsETd6xdmyXFInTmx5Fh1L8DuOXVBKsDQX5T7PyZg4jNZBi
YbCHGvqmNCLThIjBwv1YLVvQJLgMSTTFGeekfgbGRSLmMpEtJYUN+uNsPh6mWz6Q
sbhwNDWC4cMhh0cjtIdoT2anJXq60bK8iVQoqqAyGU5O4C8meZ9wFc5A5ITLW9Hu
3JSbs1GpiiWoOdD+0OgBORKrjQRzLclmnTwzYLqaHSSteom0rd2lbzX8laHe8EZl
liiyYhGzPAu/3ISUvWdMd4gz8Re+/MaO0dh7gNgDdp7/rptYKEIc428gxMaUHemX
rx0p/ONuEH42RLFChXD0w2C/b5+Ajec87+knt/Z3IDlHVa27a2Hx+isJ7FxF9OI7
/yrsvgC5VsYgd/zprfxYKzqpppsprbCUjcaxCnab6HrdQ0vbeeBH6/G7bfP7UK3k
ntr/TEt2Zo0ldZMHehZqpNEWeQpVHyHCqH2qLY8HkE3RmlBIHh/unk5JS3VzLQgb
yrJE8dStCCQuiX207NfY+ndWQGrFaOrtGO5tIeq9NmElPUHDfUF308mEFnfOJF4v
xDQBCalxImPgGfabirxVslmdGQnHhjTWpNoCeqZRut5DdWXlq28AXnj/7nFcW+Yp
9uni372gdKxOAWNXPdQZXvQc3loxvWb3fthjS/4vSCRsaDM+JBOdx59kzQMMSbRi
33QxGrC49GeX9UAua8LkHqgAUxLO4pfXZyJbvV1ElnrwA+mcT+9k+V5kzKAfrv7r
ASpbK9v8mIaIZeyROv4kkGJTvloG0RdYtI+kNxyTBCK+CQuFDvYqqxxcF3ylXxMV
Q4o3Gw1kiz8p3gwVdYlrhl2Jab1Cu3Ze+SzhlDCdJpKfZPKcbMAsBwL1L3foOUA0
6OEgL2y++dMSwJk72fRpi1plDlO7iTdj2snszBnQv2Pryi4HtoTc53W22Kkdn+Z/
BP8JhowLg6W5GhJ1ycrkDVo5jNjK1V5X2A0rYQUUG10KpTHYg56KVNiI748NbvpG
9DAxQuz7tS78fXNcSZisZy6rigrPn/yK+LWSW5DW4X0v5N9wd0v1PHCEKtD16Zt7
ChQSrazhV2BQkLLGspzwHCcics8EXOi4AiPfhiaw1D9/vfsf901UqMZ6/Ke/Vg2A
y2nfQKJF8DI48+Q/ncVFLjA2gDHJUE+BA8MHVAZ7GbGAU6ErdI0MeFAfwhsk3tOu
2oEXnMfFhnutpkeSA7X84uavJ4+m2d2B+felZiV36WL8KppsbokPAtlJFJevnADA
lC+JYEfFF9F8mhqda1apEHwkltGqUsuNwgokokrSLZ1c5TutoJmve7ALM3hnwip9
doF2EZUYODv3rA90ADSTqI4akjgWzbPfN2QcrjDqjV+VNBVErAnpnaIBf05zUpQg
zTQUrwhZlpYQr+3Ie/jXh424Qk44Tpbp4yqT6iJ1cXjaqlI5/xqqMTw/o3ePGeJn
VSXPB7HeJXQ4lu+WdIjEg4yBHGRdQrxH/3dxvmcFrpK9bsvCJgkHda5uynPmESdA
9HnVTGWTgxZD+tSCpyIjRZTA2TtyeM8n9nNPDAWOcO+onNbi7BkCniBWWlHn32Ss
fyyWOLYByyU93Jndx90DXua6u8FpXMhuJQo6fqlgSk22lX9kvd4DgCjTfi0lCaJy
S5Ex1ZJEgAiwuc/h4vnAAir11SXNjaZ0TLTGLDkC2uQs9IwwEZvPdn5iZgFVC3CV
vWltyB+SnB5JLFG/T3v7LnOCF/Jlyk034ZlDYeRkpX1G8qeZybj7BGrtgYYNzor8
aRpQ79cTaEL4QrWjxilYfSvmKILcHGYnv3ZfUhGED3+jmJjyiXGMcrfef1TUvTjb
4HOzutBWyHxMnqd40CJLMWZiRxVgeJRbPvmFjWxfZwqM76vnv74dRnjkGz4SUBHy
prPArNEHLifsirSFaFB8Hv12WMno1JdnYx1E6Xe+BklJ2Syocuzb0YNhReSVHYla
Cxf9uZV8TD+M+pKgJidvF3A0ZG6wG9gFOtZEEebBZ4brSMTfT7d4aLnKiesTl0Kg
SOGupfUk2siVjTafW98oS/yic4/l680eWPoaFbj/qEwc0f1Ox8zLQaxx/HqkKSe6
o0e9FxuKQIRN+SWUaAWy1G0Hn9ITjs8ICuE9047PHtuaoTueDQBtbG0Vz3CBtu6T
nTY8i2nOjmrJsN8Nlh6mj8JkZVmzB1UqShCknjx767KCicEMZGm7cJFr7yZzroPX
gicNmDzEa+pczuMwrWS3j2Az51wIcdIZX8GSYLMRqkGs7gE4YN0Wr5BJESDhlFZ3
f5egBuL6/2d1NG640l4ALxiORO1pF+rQ6MM8rstpA4/UUttx/IZllGuHej3cU26E
kXkWR7bPiLa3pSv20Qeq0sHCbdgH4tkOSnsbQ4oJEPL7CwQRbewFQP0T49eydLUI
dqzNskMlAs2nVRrdE+P3HFjR77WG2LNL+U5GEmksdvK27xxXm1wqyIyuQXxH2VJQ
nsYPYJ5czBqyS8fTbSog0aHqgoDXy1BA8KOvLoPEP6vijymMqOD+1juoi7pfogj6
/vIT/CEwqrRQ9f4nYdVwZd/VhYqGJXfWTs/mYFp/3e/+RRlSu5LDDWg2ReqIsZBL
BN0BxKTpnA5LTrUVUaNzZnM3iYBiHSYs+NxSSbvCc3QiS/2uBPBLTlGUBpWKYf1f
VwJaIWd8WCUi4Xdhx1P9TKP9atkJernqF0xfwWk4ETCQ0/ZnfQ1TeL0xGi0bFjRe
i/YfV38VkGbfsZoFX32smNiC4FF3DsQjqXoptfcJjgyr2vIntM1s2Acxogs7/hWE
mhG0BJBkc5EL2iRpQj7OqlOgZlF4K3uyOVWy5oLIxWi2kv2/Gy6zjrTRG8+mIBD3
WrhOJQ7yp0Qfl01cQB482GqXeROlqK55LsVbHBZn5daJXbeKoZKJQcZRhLtJ4rA2
nGwyQrpznuIAZYKTpk/PmCIAm7KsADWTM5Z5RcWjSTYAhamP7HIM0o5YNUxKJFMk
fsNahIkuDrmZA+6cg6/nDCPvVVxzFOgYVPYoNC8DLKQqyZBfIyQYE2L4L4HYiC3d
/IgSvCm0Z7b09hbsD/nDnvu+8gTF5BnnFNJ6Xu0eoFt3QVQ6WcNZasoUtajuJj3L
r6al17dVpULt4tkluEdk4wEtyO+wv/zncH88Z+8R88qP2OL3yBOFO0ys6AK5Gij9
eOLh4vVbLDaqf9Sv9vjy0/1Kg+OrGZtM3sN62qRJ3Xo+YwF3EXLgNYKMdnmD319O
hV9Q/Y3dd94m2mMzzcjADOcGkoTcQJHhyGKaRW4XPYkY687EfmXvxDTHsou/xFRa
vOFxKZnOhx8U4jaw17eHxSDA0vQ+UChxgIaj7ptcZJfmqHQbEPWQDcNOTuncl0gd
5C9UZ3ggbY+uC4h6DtUwMSGjOBmpTDeF7rGuRuuFdQD/KojFiAlZjtABQjp7VMmq
43JtepRum4njerWolvSAsp7fFH656yp083pOCqbfo6FRMXJSNAEeUYEoNRL07eOd
LvmyHhHLAdKbjLA+aQvpmBfjnY2Gqfp9qPkUs8umOdqa4PdXAYvX2lPXMvMvK4fH
E5xraXkvdZQkM8okK3x8ZDJm3x0IhPpjmJq3xntW9BQIHn/dWpcuX1hQ8rbBmM9A
iQcJ92C07A4Dw6hC4v4z5S4JzrS4ekwHeq4GrwrDrbzrAsYBq8ThZK9cJgX9bMRb
1oOB6cswnVBkhkt7QGx7arYW7ld8arIi9O0Axyv5inckZUs7BuPIr/wbPhy5i9Pk
rZiSOgJR16RhyH2K5UIOubfI+6dLL8DkdSh74p0Nan9Su0KZ6DMbobGT0nc1VinN
nPX8aj79RDCC6xoWkk0HM0NTyA3uPWkNjHcNjhsj4WjXl+sSClKVZjgUS+dc0rjy
RKCRnT4ERv7HLv3mTgdH6jGw73nYMh7CmTchQPMTu/hkFYJ1mG9/CRy7KKHdXYub
2d3Ebk0ncFSdStjNBygxFpmcglK7nbpbZy7lUDtxDYBAg7aDhbiNjpiwQ6+gA2g7
7yV7oKYI2TxlMQVmO7gkK+cT5sdxStrDymksMLcz9vkYqZB5Vm2zxSm6jUgl0x3c
X5e6vpu+1wnNEZdp519+dmYEkNklCduklFQsmZ2Gnp3ZEhVkwEUbhB6cEMlzh7Ds
kmq2FYFyO82N+5+YwJRbWajpPm1/GfU2heSxoWBvrhEnGp2E6KD6fQSrSNYU+y1m
tOpygVhN7U69HhIYYgk/nbMdyrc5tc396nFGvDe3gb4OiKmjowzFoAZ7FFYuOB9H
yG8nkdFowVs2lxpO8Ws6J1LXOHDNzOus95V+wD0zhJvqGSJ/G0Q7LuvbefNqMBaC
MPtg8xfzgd6K2mUkRNVbP3tS+VWfWA1ItqRuSvnx6Ld5LGa/SMv/CQh3+65cK3iA
APTGpa7uMNIQOBObvrfjKiElLp/6bxdPJWPq3DYxkjvrkfHHsnW6rME7E1WT2On0
KeuuJX5+2QH9of77pxCfKsvQC8yjxg75mY+6eKsJln+Hof3kNeKPcdpkXHgi3/k4
l4UpQ1EycmEfwVYw+Gj9M7xFDeTy9x4qqgSyzTXSGxB6pL91wQqzE1B043bInp2b
/wSS2LI+WAfrw0VLgu4eH9MaJ6WKyD9a3YPq5D3lSvLDBbWJ+pshL5F/G2alX8o+
VqjO3DE1ehf2a8oOAc+WlNxoZwCPeQeew+YZ4pAYuWRO+0kXENqxKOrd2hPU4OpN
SksHND8GfrC/dthCSRRAgKftPqRMfLNli8lSEOJLF3mLHKCEIkpX5H66EuGHyU8d
aKNAuAYIt4O4V30CNmOBMqrXMFpCKnf9qEH8hnnknOlysw2yXBEUFoeojPQ87hpG
4xat5t2QIQAdIJofGMw0QJF4jUOV5A92eI0cQZZiH4upq/XShAmATSCWeXUcTTo2
Uw1N3n6lMkjsRSocFDtfvjogGI3lMS7rKuiYB7vwNVb3iIsbQIyVvVuIiqe/EPlZ
doUlPe0JvDg/KlGQqu1995dnqftX18TP46N5ASoY9R3SoM/c5g5U5aDZFWuWw4H3
3t95iwPsKtuLh/lUPPowlK63lwjN4AIiM22W3c48DuPnCfYJLDYF22MtRyBtcA1r
nZOfhjjBkPRHUaKz/B0ZXyhSwdGQJTFEBG5KyApz2KmXSd16dxvGRKT+R9gHaSjn
rRdnGHPGY6h2ngCI5M4wLBhOEZnqeq3lIcDUw5OwMsjGU6QpQ2/pWTkixELsofql
O9+ZI96E1Y7/HtfT43JgEAX9VF12imBrDj8HZFmfWhVvnCiscR/EmOLY+mUBWlc0
cWKcKdacm6WCnweI71mqlH/M4ZHTxfgoDY6HSaIxX4kdT1i36AsKADh8oJMbG3sY
kdYlYotEepd5qCvgCO7LAZGplnHkof9krqnph0V9ANFirSmUq+u04Y2GbP5m1gRM
+H5Ij/yqv/pWkSs9JmqbIL00GQo31HahGapDvP3j88UTMKJQtyaDWmEt2XFKRw9/
1j0c3619A430HhAPaklLE/tr2VM2qdY4S83SGdjGYKngGrRfUqsUH91Mkvo/REgj
rz5jSQCm+CUuoTuANs+vSkyUCrj5bhRhpbZieTgi4dhaDlIUTqt7lkO88EB+MSUd
BXU7zFcW7L9UNL/3mWOrQ2gAsPLo1CCdWAS/qhW6gQjUrGZtp9wDn6Ax/pmE3aqO
O5E5qkC8/62ILM/npA0omIczMRg6gO9vX1gzgzvOcJxv1qEkpYMkNxvAmFUsi36T
tB3qJw+WNgxIGaEzgbTUKGjaoS5bBsTokCFQW8wRBiWdUR5iV0ecLY9PhtR+0TwU
HDSpMRNrWxuwB69hj9Fpf0Jkgfoc5RVgQRbllv1kE5i8H2BvHUov5B2YBV5eXLEZ
61KMScqi4n7K3GPyYVTQCfF9aQgRX4sFYlRKfdY9I3mDDCx3+mNtJ1K/DyOAMiHB
LQUGCkGOBnNb8sPPtzA3P+ZzznLOi4lPXM/JsUZ35QBpcjxet5mgBXxtWge4bPLv
wV3E6Y1MB5mZZFpIBoMn/SbG4se9AO5t8/xE+VHPQeWW02wiQkmqspek9DPJZT2U
gR8S5/nPoCdEeFJfkeIfhoru48rqyqraHfHOWnyaMnJ3r1d4iHRSnr/nyYENuoKf
aCENaynzQZ3Qxv3MHORqC+SONImJgKxlR9i1gm3UhZ5NeUULvBvjkNQiC0Uv0vdy
jkOmyv1p5tcaZzBT9Rt3Gk62EJQLi0Bg/OxGKex5CJsr0YBbKVwAbV8nZBk4vtu8
GbTS8oy9WU25YeTBx5b2aC7tDGCIHKWEmxEm4xN7J1/fBn4EMCfDbiIPMly+X4m5
diB7rgJCp7CzVjJMQbeihYHZurCwMsgS9SueEb7bEde/hTMPn3owvBg6B1eEmAbf
PbzETu63g9I9wbd2lu7TKsG/4PEsH23kmsEjXVOVFXL+wnKXMDuBA0B2KmIQKuCq
6b9yEaCCdz4iCwslNyJ2VHQ6yOKVVtrrBmvejJIZADwH0dmbA/ygxiKdwLFNi0Lq
7G6hVnTDwHrw98kVEo9Z5P9GjHr7aHep2yRUcRK9FT61qnzrnmtIjpPriVJJfoYl
2BKHOBSF1iUinfaiXpPSIrTOAmzA7X9NA9Qf2a7zwJQG+TNCYsvbmWw8X60gVm3L
FNISkPRSh8fwQ2aj/Hj7Vox0/X+Tyvu1AA9pXv47X61CvCasYGfC37UdEBE5ZNJC
OIpi6Yjmex/CgtskkEWv7HrxSUnF6gG+23kTkAFLx9NmpRoq1kQhfk10mSjFFL19
YBwFMCKsJ8fB/11c+0jPsn18ne7mrfqbfJRL6WePp/Fqqu19k3p7SaKLJo1J/yar
Yjxmwku/kQeuhPhiyURzk9vNmc6eR0UA+GxURcY/fRGY+D9dEK2PRt5UOL45s1+0
XK0D1mZYz0jNOKzAGF3cDReWgZ1bExdKdQYG2JohNc02Mjmz9tVBd5sIPZ0i7FIn
vMNCDP9d4tpeSMJxDNXn6J2szy6jqIqOwhuUc0SgCQXwmNc74SjVlIVrdPnKbrB8
gxCztW0jlm9+1AHn7hLVy8Il0hfFKCb7snYsKCRDHJUKC9HHO6R15tvUmZsnsONH
2ESEc+JyVyKUuV74BBNGjmkWidSgT36p2x8PyjU5+ch/GHLeHThXFquCLSHJXM6q
KtCjz19WaE0r3rOnLu2B97+nFchzsiVs9QsJR6gysmdOExdGb9PRQTEl2RInoeG/
3pXAqRRZlT7jhUVGbg6MFJq2XSUMIDTjvL1vTuO/OyeKW3BLpafhHRCVclGwF48V
PRfQveEHjJ0HSPrOi5CcgjDWXg9oafnfwqPZIhCUbB+yViN/q8ULL9cX/eTy/O0i
bnFn/s5X1G44tfldcZfS8vRCVx+kE0+9V8K5Bsrk2QcTEqW/1+1Sh0WwHaapfP23
2N8brWYCxtn5C8/eF4HeZzAgbiIv1Qy/42C2keSgy2koJgtXNFwmhjLs9h42p+Eb
5y0KB+MnIz+AQrVsYmQEBcphUnSfB07gaoYGhfutwyJ/gQWAhPRnPN/UHQY3Xs/u
yDKnU5zmi9lvhLG8YR8rYM0DrLrvS6+Jq7nphpqQyljYWrAJ6ppE4L0AjmdGiWVf
C7kx3CEejAk9+bWXtzwaiM+f9QXuZlGkETwN+eu+NRAMFQgcl1QWdO1uMpbOK5jc
k2Xml7UOxc990QI0ijxQ0XiXzKYGXAyAnFfw6F1ZqGNwfSn2+sXiMtpdAm3K9LQ2
rEzTjr4vS1sI9C3mOg6VZ+zbOhz5tpqao2+g6JUA0FftiGYCuSu3LgySGjghkyMG
5bav9Khm0EJFthtQzkd/95tDS1DUcF25MXNruR2ZseDFbamTuBXHPfpvgYFPb9ao
ywgNJS4Ij838BUn5t1y+i9X2Tc7K2+MRDJpTNQM4PptPBNsy7QwtpaShp8k7gxZf
PSBYa6jwmO/xiV2cA4gxtyvON/Ias2BUpEPajV0aUjL2RMcasqKYuXJjHgq9KmOF
+zTC54PS9wZ7lXWprPZ8Rmm9dY1BVUcxTfcayVfmeGGUEr3sim1zs3tyO5fz4OZA
pmD1PY+KPrZgG+nDCf6kRCRIHJ6cEl0e3qIMY+ifuMNhKOCum1aT3qq/OVQvx9oz
KfYbKBtI5Rm9ZJn5q8EtZWMRuNl7w+VbH9FGtzVpLKBmPwIs1DH+tCQ+LZwfCdwC
AR4nEPLcHzuzQ8jKqz1eEDOg0HOb+I688vy/jWHWFysENwbN4U+NZ7Rkfis5plh6
O1IaT4HDUXjIntyD2EKLucL8x0BNdGgGNc7HZPOwbgXIZBYCa3ItOVyuWhdbuvUQ
T97JZkx81D4EYAnGDgUQMZDfkJKL4+TFTbtCgXpuIvLpNEXM8iLvIopg6Eiccvkl
7bpTwUD16hxX+RoD72nExOAd5lCAWHKjS4TZqgbs7w945s7KbW1fLxiFu7CBoPe9
KpaEhkAomvwlroRlm7KlqLV0fZNkFLk/S7kYpFHjyMfli+mCMdVMFDaDTh1HMPYl
4UEX7Aki884EauE5DeoSDrgijanOeHhXb0mZ9sPzns4ApYC60eaZkEd33g+OrpAD
2WD1sCHSAH44YoXaAzz0OyJdar/yCtGCZ0jWFHw0TrkeDNMIkoFZCAKyuH8DcbUn
FiAvoBmpx7GhZnlHMGU6QYAWJpu/nzxb+WZjo8+7Myrn8cALNUDpRXj20G1lHABT
FLByarwoSFtpPCDgdifSeW+OHbIo+63/0IOb9Qvkg+sCHL5DwZ2LNmazjRtMU4eQ
XSlzxJX0hq/WCcQbVW2fwqDpKRDlyHJxgJiyuUkPD19CwEsPDZUsU/cLRKgb/j/i
qAmFD2MxP4suFnf3BZ3xQGFzpj/JT3ZsEWeVYWntineqXpvBXOFdYOGGp6NfFuLk
eApgItitDEB8Zh8Q6d88fUu67XUnQspDNuzwamqbtVri9DWrAt9orjQlcHK/LHR6
poFrG1/qsQgaolqYXStw62AkxN/OKtYktZltoxjJsMMYjfjVX+nMMNRbByUVFrVg
tLWVGcp9iN5u3e2YwAyNWQdIpVt1pd6AZu1UpsBijHDAgENOvW5Ct5WzhsA7Mmtc
yZ00cI3l3b2tql3zjEuasRr/b2g1446knd9INScxszgqD1xXJ2uh0oN4txisjA99
/OB1L2vmxguEE/deMaCme9tMLo6eis3fPKavgftczl8CF31nmykHLz3AvZmPBihE
ozz7lTbOYloo2P94UTzTfUSJHjQEsoqtNDSHvlhYYjAtUg8FBU7wgNd/KMTkiPGt
9+xTcvOZa37htzWyvM+sDDXLryZ7j2QyX1MHt4dU6NXAisMbVeI9oAXEz6bqATEm
GezZD8RK9HqAqaEalSXogiRboGNG8cB0oZ4mDBbJI9cIc3cxgPwdqN5cZf5kfikI
FoFns0jCeaHt9sJMrgQO/dYGsZ2twbRVNks2Hn55t8evjGvbAKbXypUMLKNTbYuY
Gms8FSF8IPv2GKJI2l0Bj0z6il7Sxzd1zFAHVTLQhoPYTemeBkN183DUc5Fr0sY4
UegzwriBx/9T3X/wtKCTZZijMo8cvWSv3BPdxXG4X2HiXr3YBF9Yu5xJ2B05/zGQ
eeFSKwR/nvmOSYtS/m2bxmPsbp2t2h930JL03/3kA9F0xk8h3aBto5qRqqPoyhJI
3N+wWKNTfBje+ofGyguM3bF+105Vizb8huXed6YxgkV3gfH2nMgCyuuWlrkWrvww
DPU2rTbP+ImvY9/MkWgbHoGA0tFIv+mC9yc4moBguQ7MMxDZCcKUp7Okgs6fxM/l
2t291IopQqdwuUQTy1QdT56GGGGUINkWqYVdNWDHSNzBnkLwKrjgecd8BAzFJFG6
XxKn/JL91k4vP9Og0/5jYdNMcg8hTZoHtzp024HlWmKd4c7QotkDlSKKIRLyPwGx
ie9XKO033XEsPOE3FFDiP2zXe+UokplMGqCBJvstdXawHsKcMSXIxY8tvF/LkORr
rkZclhy6CNLl1Pm/Vhxg2zBDS6Y8lotvNmHFd5iAD2j9gQ1K+wOfg3a2PQDxjnlj
lrmfadKkGsT5g7Dsi9+zNqTJG6TDLU9fiQ0dXbhN7j11jyDo5xCQXiqvoAC+tMcv
Rs4I2/3NPdIBhFLStS2ngSzRFwxDkq+Zmi83ZT7v2ZdBralEu+fe8qA7A1MtRumK
Lybu9MtWvWnrnAkuoT7IAs3MvzFrdBWkR/sRfBHZ/E0HrLAGrogfEl7FH/qFatUT
gg3V4j7xWEQEYWf7ES9FBWE+5XShdqB9LZcjkzZuA8CsPatYLU0LFgdcbprw07e7
2WU39gLjtsOB/ziey3Tj6aPx2pB0zu2xVMrnD7dPBrChqB0n8Mtu/p8f0yA3XJuB
edzrHdOh5KF2uvCaOsEl3Pp0a7mVFTi5huR21O9ZbJ5cPKNNPejOhd8du2nHBq+h
lS2REIdK7c2BsKOCozEiSaWmQ3huO37548Bm7J8fkIeCoTarNjbd0dUh/rdEx8bO
3XmZRmlRCbFqUjylw4ASXvRcMuucDC9mhB67sEk/IvnUhRm1xcRZB8kGKK2hImLI
amVZ6N0l8nY9A9vtCegVFi2hXXPsr9r9vUJvdAFvrsxBFIu/AdOft80TZajZ4Sci
8e+CJ1/NGgvS2C8UXnzvdyZ7dG8DJx7uokxWT56UX69a7CjGLExouroF1mK6Krhp
2V4SRLwDemY50eXPIha4J9CZWI7f0EANx7VmYSVWxl/dfvfoAQPxJgTQ1hRkYpQT
uVBzWe55mBHIh4vJ92sGkDyphh7G2No6kuJqiZO2sTAaqH9H3Z0noX46dh5XaOHY
TkWQzRoGhUUDN3N3UNHAYdGFIAgjugINLDnek0VTfYrcCOLP8kHxF0M6mmEmqeRY
tCPgorgeb+yN7odiRQX2wcy9eUdMtoaHrypaIrev/ptE8T0gHLPexK7U53LBHApW
mv96KGKJjeDZi9P9uTRYi9qtEZI5QA77AdLVhgSrACpsWkAm6L/ChzLD4BhKhp9y
xKHgKhr9RkkqOAe/D9tyhsfS8RIUmRdMutYBAc31lXVzv52lUjL4gWT5u80suWr6
i9ELPe/BSN99oT+CykHt7dS13PohO9kxAdz6vgSeJflEmZqwc0S2+ECs25pwU0fc
/wp1LdG4oeecL9XMfIDiatL+RpJJw0TEX8hVK36a+nggxeEl7DdLrLtnBqs+vUDn
7ooTlHGvVWnYqOV+vFa+VW0cY43bYjDC1mAXq+L6Z/sMMt6iev8Dj1pxYqGe3eWF
kzU4XKIF75hikq4KLKXqwP5GT1V63Fw+FnptY7LODHixpXN4aYJzsMtFkKVMCS9A
Y6uOER56XOnynQKqttPTLkM0zVztvo1AyYvbUPEC2SazAPrPmSpBFQ2ZNHla3vDy
AkGcIq6F4gWT5+9t6jkdpqJBPVdzLEiuz0DUgqvOTl5dNEYwvMrU+ZjZTGb7Je+g
IzLI2E+S3X4pMD8iO/2JdRTw7JCYy5ATu+lTqtV3QtJpuiYXF+kj7KQs4Y5Wlsz4
PDFNT3H+HU/pb5W6sBWc6abKQgudDclYG/Z9LGLrMZKdrMGWQwO2kf1KjHsu8hm1
25J6vaTp4AFLpEJgtMCDuxO3uVJPAUeQevOFt7znJMSjjByAvQ4lfxGO3ct97joC
Ke9NvoBq+Rql4lpxzRlxPkX/oqAuYz2+AesnFzf+AeitlOHB7dwKpf+dza8hkADI
CMGWgx0PVDXDBozIpTCPD+nTsEvnEPUeABR9RWv8+PHyH+Zyqrayz4x+i1IrYl79
SpJqXa4EYuFKmRraYNESex1BsjTBF3ng/HhauiyueTZKx3ozwlAa0XBRLpkKaRUX
xbHM7szueBg98XMIuwV8DtvGt7JyCnAjOjcP9emJetVXFMyGtXKvqLD2QkS4BgnW
cclLRO7i4DqEMVQ5FrqdIsIa5gP17PtYF99okpJwb6aJ/6IfdiVhQKJrTVx9vUkw
zv2O2xyeQ2Dn3TaYWwZn0hGmiPJPlcNnOT+eLxJYsXrGciccwdGmxRNxk7Ea3C4v
fL7Gnn1E9VYNYRTqj5Zi17CyiOSpEM9YqfUdxSacXYr1wNOGkgLiWvULybZ8K2ZI
zIf/oCjFN5C8DHsMx+yv4yvfjsuQl6TIDeNywFrLZhRQSitK4MPpOhNe0uUce88b
brIxioxSUnNv+uf+k8Zx9GPZOhXgbTH+/tjFk1bCjhX16Xyzr/fAddX2U/T13YbQ
wNoN62RgyoUm7YDFlQKb7x0ffim4f1wc3Xt7IOh4KtybaPf7swx7UTn251kyqWY5
uC8jBn+aerBxnsNWTtNw5n6ilzynYu0LNJSvypAJdaJ+xsQSJE3ncCGAJHqCVfrm
`pragma protect end_protected
