// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:07 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SDLOyKb7p33AooomiuqgGLIFf0hLGg5ZLRyOyrxoLIJQELAgNHG7mFckICukNBAy
V501+X4DbVmt8I3iUkLSF5O/G4vBKoS8gJ2eW0uPzNYELvcbdB8bO8AAJywoaQD6
Y1zP3PE4c7mpNmk4ieF4HoEQ2nBA8E2zLmNGGI0ALUM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
ycYTnCopn7VMnRWlXyvFX3T1K6CSbprFTNgUafO/c+TPXbIU7H7R7nkaQvAL8SOg
QOwJ7cGA6sE7VGYl1zXhTmnUi2UcsvM60/rYpqaLIIoFLn4J+fvlcYWzZysPFsOe
wS3DAzCLqe3heRwcqLZy3nhMGL5It5mAZzNoEXdNCX775iwZIxlDgNeZ7pnSX4bD
g80sLsXKTYlTW8WEXAmXOXZwbpsSRKVjSJO5Wiy7zwv0in6k5ORdL7utSZIZ5JIr
TtF4Xf9DORVsF+yKQfGgzBoXESaXKy3tPmcb/MPPDJLF8itZqGLPuianrDaAxR8p
DwR6qYrM+kb+lih6JaxRaNN9wZfBYW+Zi2thg4Gu2Xcd+6c2Murbgfky7ADmDMhc
v07ZkRhYF8G0KCKceOUj3juAb6KmaWHfxi/P05Loq8mIYytIUcQy7+D4AbLa5Lzg
ENkzPdh6nUqny8q1iifg644aT5R0Sg2N4JEQe4EsbSpRVJhpWKoJBVBu1SrSZhiL
rkErxZFustRxBh8g/uZRac7yzqbKzXeOtY8ubE6kcWvezduggGpoOZN/XZLEQosj
iJJRrQYt/4nsfxbCaBnY21W/JrIrHEJgcmSL188o37jQaJy3BjyoJW2vfkbX9d9e
pJfcOJAiQ16jYgntAfxBRyzQXW85U164QZ8kY6Vck+2itVpVBzWzrWOpqwqisohJ
jO9yUrER7X4MCaM0a0RbS/OHN2Hcw91zqDRmETWVKXybkXqmWlhCxC7to1w8U7oS
iHx1K8o8V3yXO5X/X0l8p6aW1YG65Mu/7C5jAE9jZnBTDQB5/DEDZwOBJd/JWUMy
vnOk0CizdDWGV3sVClBrLXA9xo063zDiZqq3JTfmhl/Fc1p2wuHntfLkrA52Cwqw
JhYgirIEftiW4q0woaXclHw4Z54mtZOcEJ3Pbtyv3e/Bx8E0F3Xt3esdIMcRKFBI
n8xiaEwNVjrhewpxeRblHCJi3vid3cl/vKu1SkF52AkjIqBlE/F8ZQbl1tROWzSC
OrQgj/MtClLzL3rF0u/qH2DpeDb7zhaC+edJpt24iyl67WnHo+E25+rUpsiTmwmX
7uB0lnGH1bokVFGc7MWRsS5j2o2u0zyIAqS+z9kZIfcSmgMCog/fCJo1ufZrvLme
diANtfuAbSg7j5K+gUbpbhr5zZ77o2jrN2lxcEbIyK54+C0WJtiIKfMbQx+TiFAv
X9D4bTyL+/NbK18mY8UtGLKyYIoCQR3EJBWHebmbOHmhd2bRzuxT5psTihssbniZ
GNhGOvbiu6ZhkzEUbsNzpLvKJgSrrbOVX3G8Y6Vlt6hMREaHtplW/z2eiHVkaZA/
yRnux73Ln6gMUt0sE+z2kCzVR1LbAWVnALunfwGvn26vWQHtHn76mGFOcQGU6CYf
Uh7ymuskje08S8QFcCQMVtzBWxgvy07LszRZWVTBtlyA8B756JkxhhrZF0NHHP0N
QzjuSlgkGyRfum9UR2mfniEqSNeokTcvt+Ba69oYV2zb2ISzntW4su//9tBZo/6+
Ib1R4Lg4IYC+HGwMxlByPMl10emGZrSfxnAfC0o+UxA+7j+yHo7F7mqLjpgl4amE
7o4U8isg9yueDslNTihzFKJ1aAxGAId+UL4haAgdn44rnXyu9kAKEuc6WFgk4S7q
+7Sjm8cpxsVZD6AJUfR3YHcIalYU63xmt9twcjxyYRxF9eYnorDCWh0Jir7k0TJm
aoVi0GfJ5eByzAjSfWTBNEtNg0jhMr5tTLuUWOTZ6ckLSry9LN6Kg6piPFRsq6Vt
dLuYkVvDJN6RPtlBVIUGGC+7H1YxSx78irr94Zg/v0eCs2GiAZyNwdkMmND49m1I
t4afeRySjIjZz7ZQja6svHGOp1lCQ6Zu1fkxPZQJAmMnzfaxXlE2gSD16OsvLzmN
LNs4iIwa1Jn1ay4C+N6AYAxo5tzfxataDbi67NG6J5vaf3B1MlB1RR4L0pcukxeS
nwqeSsvRR6M+0znWLT074qr44ee4t45FArc3qQyRd1Ftgr5JAUJMqvMene5Gvpc2
T9gI9RmYau/VgR6fcjorFe7w/E5S+26KCj0qn7IOuWWMdsZa7QDmEZ++VYS44l9D
zfTPuc2kgwJ4uGSR5N6GOiS2WJyJOvS93B1JnkraTTJjFYCLDCP2QdVCEvqrCTxv
f5ay6F7HZOEjKXU3ByUWa2oSHYtxhlX3HKoOea46V7Nr5ALE5bKf61vEzD+dfaOS
gGrQfk2T23to2+kXrm7QkUd1BQZT5WibNWfay56l0pAC1EsYzU1PvUkfyAJRdbkF
JMYHE0fcUZS+f/e6zMCN5jCM0dpZARTIrJObhX6JVhnMzmUlXwYMaV+JSmzJd+KW
zCrTaZaibA73WZmhAOn1zNZeKTi1k0JS+/+sL3GIYBZcftSp/pZJzMs0/XOimeb1
XukiVgFCYzBmqaXFexkzfWqAmxo8k+oO89oKPdl0vvNg7Ncjp8KJK1Bs8sVCLq62
RiO4yTNpf6HMzuK2HIWfGqP48YTBBd2sMouI4NzIsif24kuFI7LSq0Vg1KVsMc9l
LEysikHtGox51xdDB/vTh0QpmVhymlr1c5vggK4PtgPWDQEPLLUGHFGmSdUR6bWo
jeTemDaRy2wvfmn3IOBEUSiy9+hOj9vJOGVZa4EdH46IIBH+Pg2aJ6EUxR+BqJoZ
cxNtc9QvBVaHRZeW35hwXmO5KB/fwa4AcSIvatOG8uBJK9CBMoM++9gh7eBBAl3q
99RXHhEYqic1tP0ColmavKRL9hE8/Mt/Z1VvHTH/vAyyojiMvCmf590EUYxCnErS
OzLMFzFPT5YuLgYUCjbxOXKj0dHkvF6QgAkOMuaiFNfT0y06Qvihcgot5ZujHa4V
p9HrTZ9NB8/UdyqIOKP42WuV/eJF63xXhIP6OUvWX35aFRhwxzooCy0P2zAoVqYY
h7s72iBkKDfwX3AD9eYuIJz4WpglkXASW942vxYpFzAVKrZANWJ6Zd1fM9LXS8Zi
2yEqM5dTx9pmv8g3W7spLRH6O1OcKutKwwcPz3u0hiLwxP+OvE6nAHYv3yox1BMk
RKiZ4sT/lEsIpxzohXkey/UtVFqKAY1j8OD6/q6EqRujFGsdNRvvrjO3igvBgEDa
JOymK3pZffcQcHZfWEGinDNqKEF396MwCMp5JpUPaeVqQaLNEtN7Q27KRUerlqZw
WLLbKP1ARwXcXHWsvoxwPc0a5uwkGILjQRSF/DCrvscVZzJpyWouR/HYGJQmzhm/
ZDijHqL+8vZRE2D4I07IUN5VbfpCszqvn3SvwQS6MLvYgEGxkgZvJb8V8be5paFO
Uvt4mwsph68sbTIzd+VHc/c+ujrz/eEdyTZmmmgg40CDWRusiuT6IIEcDfWqjuB7
OAGN91QrUmnkaWvVGc55YhPiq6qcg1Uz00pFgX7XcOGe49fNkGgQOByrxCuE+Tok
gYbQqPDlzfHHUFriVgcfKbdwMX/Zoc4fM/YVX4zpm/rda6SLMirIe2PAQ1SWIiw6
9Jj3/0a9t7eoCCHW9IPdPeAVFKHe6BixcN27uwLeAyBJvFk0RoqC2/xeIs5EIPz/
fPU2mJSpTTmP87qs6IiVM13HMoNYLpMDmGB7yyEZmgY4il4g2eQH7pbFavUJzrvR
G3f7ISHU4OsOURiP3OAA32oofoycXrC1ROKybtKwRw+UT3X/AGRhO/jw8E4O+TZI
cQBtVW8xLU3+UrAooXT3lRufXyVFod6qiemzVDYFzg9l5Iw66XCVXU87LIErifMI
+E7gbjI4BdsKDoXIZBZmtKGeXMuk0UMbYG5dkzMY0P+heE1MT2RMKacmWisFtIVI
U9xESnd8ArvLP3Kt6pyqq/a+YUzAWuT1ZU6VBGn4x4yF8maQcMnCaXgV/z1VDXUW
UDpM23mMfC78tgOiRHIzGWr8N75QyIUQhAeaqsUy89+xO/lwCtgihZw8SrpswzZ2
ACE5SgTcerEdUT1/RV8paspb/jba59M+zeOV56j+AG6A5VG6MUGXH3jqtUyvYMCk
ZKaE5mJdLLu+T6iNaHvwTM3bmEhHvl/NTPje58zIGJdha2UJXpwRy820H0YBCVDJ
vO2fcM/Yw3EgMosz213ZWsfSmrTl9gyDNOvfrLszKNNwgV04lmgzIjHFgS+/9DBU
8KzTBEhDLmfFNylTwesAWKM9BMVJucGSSb3BUZo3fiU96Cv0SyNlU5sQig7cLZNI
ysrpgM0zvTs9x0LpktGEPPtti3FRUEqCXm5JJvcqyxsl4L6nxFJcJLAnxZXq6Ce2
Ymcao8NfKerNvrp6CmegTDsanNIOMRNf3yxcYtR5ko4rYZSsCoSiwyaGiqYiCYzU
qN27N5eOtPzoSFp6udH8QX2iaxhkLtE3QJVwXvoN2bwyNgZHBK1Jd4X9wlI3Uz8Y
QU+Qhc95UOm4yN2EqMRH2Z6buuv5JKDLddfic1HLhHCrP/MK91E2gGpKMnBIrIo5
J5VzS08IjRk5e9qD8X3A5r86yhZyeuJLApa0KLzcQJLWjup7OCI46gc0/ufbFO5R
Ak38j1jGo4NMif3l3hC1cdRYCMjwYC/ixBbezCfhDR6OKavw+hDehY9UKra6NVfp
+KfFJmEN5Ho7LaWSCgBMvbAYZdVeuuICEMy09deswcP3EFyEynVN9te96l4KQL5g
g5A3G7EOJMUaTfc5zhRwog8A0zkAAifyIzWKoctRVPR7nabwefvyaS5vVBiGl2Rs
UWUnb3hlzeUBHvEO8TU+Y2YLq7guApa90AMUbUbqqaC02cBS7bOh9c2ad8na+eeS
WeGUEdXM1r1LCf75X701+UZFSs0yX80ZGWAgbXjs2pFHn9pRi/8TaQdDW/2OhThT
h/dCT97gsfPKgPotYGbX3UvGWMNKlS3EmDfy2PCxUMH1mJu1oowbLCFQYzo6lN6d
vZzsg3algXHDV1xj6JRF+LwCxjSK9KIu+vQd0NwNP8yWQFmZT7NVUDW1DFHKZsl4
wyWjkrfAPdS4rSVdu+TGCGbutyKSkrTNGR3YwfFgrsvy93y2hXjhZltFnefeiMwR
pba5sDN6wbT6f+O0BR3ne8a811LzGPeDWqsQ2SrVBX17Meq/37S1z3GG7wDCieex
JN1yCqC6BpDazXmHwExFqYhQMBaRQ9whfh5HhI7KirUsFi3uwp8qg16uGsYylHai
pA+tsDBHF0ZY+HE7GjDLjxjN4OEO5DQ5lPuDVcJb3rUfKKEqgEYJhVoM9issAFau
bwNSnGtNSq2cTRpGWTU36NHs5X5hmH1L0STd8PeSeGR0PnDcRzQgCt9Q2+bKtkNH
P2stJrcVNj3Z4VoaHeI7Oyvhqrdh8EaAlodeJq1rQ/DUfCsNt9+9L1craHGuCts/
H4Uk+tIv6x+m49GTLT1jplZ8xJWNrYDGLXfipH3z7azApgnZVCYsls4wkslA4W52
7bF6WVAlJq8D6gxIOWmYQtDjbOdOlAADZotNOCq+VKvIws41t1UkgtP2DMrEXb2A
Q/pQR1dae4+rzog/ZftwQdHEZPP7EJF8a6SQgxvWq0o3RZ9nZwUtprvyeyESJsdQ
fvMZBRAjn42MCgz2+PwKd09OpG4K520WckM0j+c23rFAdKKziviPeNJsrzlbez0P
RQSyYOAXzXyd1PwextQr91Z2IwkqGx6uYngU46HI2j8d1lvM+Vqwr7AmpxL18D3s
MCYQR6e24XCHCqthADs76sFTTPVAINRqITrjKTsp5UcPx1C12Ixc1De+d0IBkaw8
hTAlHJVvmJOvPvYOaDkbQuYUMm4WxPJA9+QeRmusDA0DZRt32tqtxmgyGRoFqQt1
Zze4aCoDkftATQPnkO0B2A2cMIJSTx5F6kPfp9VNIFwmzBw+U3Lf+Y8g1H+uIXUI
/ymAeCrlWSvkWOBNrt7QVRZjM88qdPsA2PKcvd6RiJblkxbXjF1EYLhmbViu5XRS
TQ+X8SpMOZbOPQYaohaNaPcmfAttXYrV4F8NGGYd1heggy+xs31RKbS3Wjuw3SJz
6wq7NglUxG7wcFpMTqzju4ykn+18EgLmEIL3SoJnrJsu9CWajUHYK/noDAOaIc2T
eMSEVRrx/lQSj+37/ZOTWUkw4J0UmN6s3ddOuk2ASphVBDhzSrZK313Pmdb/VB9O
DEZhGpDrK84ggLgVkXz8dTFaakmUTS6ItbiJfULF6wHOs93KcU0gC4qM0ICRK385
IM5q/2/nGHtdFpWRbnZvJqHqoVbeguLk5dR3UufuhAWBKFYpsXXHPSHr081R7u9u
4FebMO3cLHX0hmZp2Ppry2sq8rwboy94BYfAky810xvBjc5mdJG/ppVGnW25//dC
HgaNmJr6I3cQ/m9hSXn4L6RNIz1oU+Kqp/yIX3bR2gTNABkEXQ3/u7EkkjCJH5RJ
z1JQ9SycLCreL/qLOUFZ8vOUo/abUTKrJA3eqgyl5Qj/Y0wyecyUFtvIVrvjhExq
z0iIs5cujloA1R8jdPU8RIS50+HOqxTYDz/0ZrxVKl1K2d3POggNt3sjo/kd+AK7
06ExXaiTrv0Y0PflpJzURFhoGp2t/zKqTBrBetLZX8iDky3k9u/JHkNHo2J/T3Bc
zNHKmR1JNMNR9CP9zM50UCbFk37xub7pIh5d4ClBSLQyUOXjD21jW6i6Pb8JE1Pw
WO8ohzi3P5cPNOerJsdahfQzKQIsB+bfByINZOHOGMRgHiU2LAIFQzG+KiwcFu8U
9+Dk/hMiFfqZNeMIKOsiLo92vqaWFJAZ/CyjzuBar9KkrD7aMNW/kQbSwJxR7eZv
jN2HpUHxY7p/Qzr59+jzXe2e4xIyK/nLl9Iy3gvYSANXMMETOgmZpFW4loU3hx2c
HYqOWuPQzYyGT5M9S+NpBBWlCxPBDXRHfGevGRoevAjlar30LTadyykIS0ATiqpX
QIqPJzdJtX7donsQ/vCTMEJYbuhMYelnxMzyNPKvaa0XpQDZmuUaW8pZ1np5xjfB
QW+4b6aD0AH+ZUfH7EJAgid3uglPA4+KByFmdLsDQNjTBIV6+d1H4zTlD1PJZe4M
22EM9lNwkY5fyh6CtEFhUQIPnjbOx73yzvtT7DZz66Cjs8ExqggN5sjjMgVBJcal
lEsz98J7Sx9OM/Zo9v++tVrS9tgDzNHHiJEjxB5Vqhj8ACfL4Ndt8Y8dwIAezYzq
fJmG7pUqG53/rkAFA14TW1aVjvJOFnhcF0xrfiPQCHoUhPEwYOAtF6jH7k6AV+ZF
Z9szXXFzC7/q70ewkp4uqhWW4G4mD1j19ABD5ERGAoLLpK4V6HMTVc6eFVb0rTn1
fzsZybBMDM3IXjKo4RKHyON/1psNktoTzktxBbC0GgBStaDe5e30lgVlM8gSIJ5r
Acji8hHG6PrWfrUciPO94q2t6tkCXAWWsWPmRzvpJNmoJEnM02wnRjtM6pKOvP1n
arJ2OxiCy9YX6KJgjWgaQFnv6O+KbxMSFPuIfNp7fFsof2LR2x1cZX9//hkcPaj3
dySi4aK56qBOZ8T9BZXhg8lVmSaoT3kwY3Ntadb1us7hkjo5rOLeywM8//LtKJJG
9E+dqHtdGYTX7rHeszr3PMj+CQ3AYlBmad9jrRlQ/SXQXeaBrpWb6NzblHp7f9UW
vDPiDUsfmFi/BKpy6wrawGuNTP/tuXNhNAbIwWd751g/p03KBN0UlfQufmYzhqiM
tN3Y7JBqgHKpBWBY4ZxOIIF/bDasL6K8yGLcuE/t5WVVwlJHsLvuvi/+BuA7r/WB
32r2gnMwq9DacQGPnq2Vs9AI+nQ4i6F3hlQJi1CJGIf2V9oYBanpAZP2KUG+Pf6t
KX4Y2mul54m9JLjV1m+2ilpJE6qerDPDkzOjsnmbEMem4bmm4FWs7rU73VNg3IPh
Ty9jPKH7dBNBE/7xiQTJAQS2asHjfow215+99x9L6FrOKY1aW1Nq83iyogl9JFWj
SUStMYycsAIfK6WR03y5bHvsmMQIc8ZNijG/pz4rV8g+0yMNJTOGu91/WkrRHcOg
sDyxK798pTh7tyBHAPRpSm5V+QIaopldbS6OJ8tQkUxBOaGhdc04MKSDYKzAe8KJ
/bFe7TNA90PMOlC13Q6Ql/lk49GUfW6AJYh/iEuhyH7RlIKeJ3PfjIN5HPd2JGE5
xL1mcxcnQEQMIqRajiuMNbYO1T9sBmQyxFe3HDmuFWE57/PHtbcTlF79aVmZ5ibu
fS/ewwoDoHCfjIoo6eBn7MBpyMZ5STZsJnunYFPXMIL7bsPcZQJCVxe3rc9EErdg
q+LSgYy0cECRY5T5WZYrSYW31bpZqHPZIbwSd5ESM3krHZtxP1x6uIOzP5/L1Bsi
IfMyjwZHaoH50v5ApYUHeTDjP6yEO1+qGR6XfM27Vyh9SgE4T+OpQpxm6pPEt4NS
5NWeCVb07FkdjTG8nDjzo5wfRRuSp/NXEX2Qorr2xVjM1LZmEpEa15NV01oQQyzy
Jl55KqPN8YXiTAwn3ZJg4w4QA59aKpKPjBMwG2RiEa1j+vUZKaV8KGGEH12lyh41
TQZEHSsOlS9wksighGVizbbvK7LzTvxLoAijVuK4pMByuDvQhqnMXMcynoS26EUB
TVt+xkzAgL7EPt7p8qthOQ96SCqKMS770OZhVhZWPYTQPiwWqDgyhEHM+WzM5WvG
lmStEcpx68zgJXL5ti6B1mZWsHuXZedhIlT5q6SG7tyBD2FL0TTfC5Nc7NmeEQ5i
9PYWGDWQpUybUu2rwHBTkomk/zNBLfu3n95JeznvXiIg6oeD1mZW8/0voyJolpgr
NsjbHrvgnGxZSpUj/yVM5E6cFxSsbE8qhpqz2d+76U3U+qfyeugVF1Td/kvQXfNG
GF7SuU7SfYFIbU7KmIfSZYF9oh322RlHjVlnLl4PlNRUOSXhR0eYwcLQOfEddOh4
jvLqrSxsj3mKyUk1jdIcriuRh/3dzH4+r0NO+uyVq7cykXrWqiWSeXN2Eg0n8Z7C
jUHZs8vRb94Vip0gh9MM5zoR9+4aTrU3g+nQM54cwTE5S62hu8qWECQ9mcGceeFP
rMx309J2jQfa1sScImH9VHyz+CS+zumHjrlD45JRwPit/bcTBjYp+Lg3yD6sIOyB
DjzhBl5U9GHlcTK0a1/PuY4oG04OpLCvIJUABgw0SjrhhM/MmJ2h6huLbF9DhMYy
N1NT0bnzFPpQ1Bk5GSV0aCRcBv4d4/NnXQULShGUZghozT7MbbsNoAgv2cifoj34
BoLy4M2p9r/O91KuvPYPjYvz/owI5VaYx6okfljHbxpYyT0oWpzfEa3VpvqydvZD
bofmfpZLRXoa1sp52T3zHIfzePDMjEuUEYboHGNkvHv3KAQwOPdQOaRlVelEy4tQ
KbZAn3r7HAWs8pJhcjnJfWBjBQWFMpIGRRCOhdpMEj2UJLmMCTf8x3A6THVs94HI
PcMjR0ldT5oa6OHoQ04JzCalqbVEDoKfrQEeRSx1x1+9iIWvuOegWlSDil02B2op
VmDH3PK4CnOZfTgP6Pe6pEnJB7d0kX4edLQ1IXRZpzyAeRFYNf14OzL19aZsgQWN
b5kvbACrCCEjAVSSDlAg/+BEWcg22DYHx+0aIaNVMW2tdaY3jYSrFxMZX4Uhq9G4
DN0uccR4AQj4dpSjVubQOjj9MHfzvalDM3mw727EH+lerhFptmMjMcE18Latz+Lq
clCwPBmM9/Vlg8K2WNF9p9Tj7MUgxFBOqwweNMzL5Y6dW1XGufe9qxZCZrtpzHbW
Dg0UakjqJ/J+8QGgFHjUzEmRQyaKwrsuGLtn4MO1lrUXruupFLMh8io3R+I29La9
WISVJu67BH9juygzbL7GrxCFb9ZtSq26jxknGZ0z3VIwbzOA4xO1yuw5V7dp5dhn
ss8f0O3Re31sPyyQRc5evwreWLcTcyjQzOBTpcUKY/YsjOygh5s+J/juurYyFBXM
RST/Jz8cumUQVKZeGK24OxJB1KTsvhLuHBUYo2QNMj8ntQnwij7Vww7Iuehf+h/v
WjNr2CjoTXVgOx3/KAfrKCzBGfTiiFh3edTP7XrlVfcnkO2TTUs8lAy/ZnTeKgJq
FElfjzRjCQf92GvzQMaUXdWuTbfTgiXffynIgMbr7Vq93jCcRcOTshpPZ9L+Rcc8
wAiUTyUi+7/oYdHVPv2MpVYlBxxg1XLKiOrEmGnLqvRCG4Q7yKe2+NABHdUL+KCT
8Qpu20nrqKAspNiIeWOrGjGis0vL/JEp4mka3eUJtuWEgWcXoJXlvzaGnIZaVWWY
M4z0x2uharMdlOqwoYWnrfb+OmUK4AdK4KOzT/fFbCUhdHoaUDTtTqhOX4xh/BeN
q+Nvuvc5eG1QC7oVVzyYh/VMzfFQijqC8H2FO72Uep1XEQOxONuacwVyOPyPggHw
wE264dhnqtFvayfmm7BE84xUzPObW6VmeMgFGkL4HI2dkegRTDA+I9j2PsYcOwHU
U6miKs+lDj8Ilf80hTPuHIiT2+CCgs81q4ejESPYRGiX1vWuKCkUOMwX4bKG/3Rf
Vsmdvqu7/oiDoGgzfeePyfdJUjNToq7ATOx9nFcl9WRzA6rBBNmgj4ncTNCtCiRx
6yVfsc0E8WIsT6A8n7DM7nORu3bcI6gSpP8h2+yRywpuOCcSsfpONKF/0DzQrD90
Vq/vhbTLTGG9ZPAIi6y1sz5tYqtw03b13DO0AdW7PRdoZ3ItZB+wDD4wFO57997u
kQYohlTxAUY0vQeUHEr7xZYNPXV/xIabipTxBPb8pvCpIFZjIY/IjE8p5+oSojV6
R9JD6Ynn1OD3xziXcRtWdrspTzER9iWVAJoClKUtd8aNqgESIxEhi/lxvjU8wNbR
8603TVkLc6I3Zp8f9qpumHsk0iO6F1XBERb6OweVTSzKr/qETe602bWBnojn9CHr
q6S8dEDRT0Du9JEmDrGNOt0bTGKNVkW88ZDYUksLS35VjcJHdkXO6Ri1k9/x/qIW
S6Dnyo/ZdVcaKEEI52OSYZasbdhHYVLfJUzF8uUZpaX3/u9IKiOaP6yIX9gKMAKb
66MPm4FmXv678ziwxvSws6FXxA7IHFmGdsZo5TxuvbZAxqODU8//ZlvKZGW5Mc1t
80RSJkMJLlJjlkEkgn5kQoRlv47LY31mB7a7JnMhgRxD9eCuj2AdHfEXLjP4rWyy
Vs6Fjf4XAIhq2CJ/pcDP5CYk9rMhaa+J/RrbfLo3Ei+eVNE6pKGAUetqo4c65zZv
E/UhqGR4PydnB0m+A5N0qi3uomFpSlXTfZmUjw57K3UyPt7emYkIWguo/mfaUIxq
Yow/UXsgSPURtPJwwQHrAVTaIImY9K0/0VIhNAsYtCjC2svDH4ziTvW4tYn2Ugcn
sMecJeayenjoGjNCpQ8qm/PB5tSeBRdTsA1gYlPl/DGmw6d5fTMMaxFR96F9LSeE
AIOxsm1PfdshbnHNmBRmeO2fiKyt5OIxtIXOy2o8DA35mhCdTwL2QAwG7SZrl6As
K6oVzMHpNn9kZjkHvL8TSlJ+mAdUGWVk5cREONYUB9KwqYyzDgok8j/i4FKfQnp7
TZK+qUulmvF0wZzrGAyWrjDIU+9urc4bvRVQLA4vhTHcABqf3e2jLJ8c/sZnTZcK
gsv/WkVQIaayCIqOH/eib7bn6my6KApyOSERdo1a2cNtpvEkdnSSDidpmyp3Xzhr
YK4ADwV8YpyLYCt+FrXDCZTnVN/MYhY6bbWI13wzRg3aZBC6ES8qO3O/QkEzbOcm
9YSKEQ4SZpIQKUxTWIONDg+64H+rz7IZMhKs32D9Y/zyAmg8rj7aoTAbmN05n5vT
lvi+5OylOdeZCTJS6fA1W6eiLnlJ0LSUrsm8hHW0+HxytuisqnHFWyRgKZOTPHIX
E4ZK6ATcYXFiJerPPYBN9Fv3PMn+zvBVWvgy+jysafRjSVmE43LxazgU+P5HUqP0
IyWITDetW887xzy9VKSN1877vUKTv160v6BE8Ebukj1aAdjk2oas3ptC4Ot5fcAB
z20qyF+gqHqnutESGVLxnF/1bsnuWMcCkQPVD1AtDk/ERNqKbXJ/iuJlcw2Y/tDX
jHD7azo+tv6+5eDZ8szEkMP7pHTLH9OZsPbs/NTeUFR4mNsamXo05WCLqRyaX4fr
OCd7BWK7N0mIBsdJk1apbIwsFO1RRAyz7TpoRZ1wg1BKmlwx11HIwFKSCnpIeapj
7e7LCvWvS3UVQTymOtDP+dWGwkl4PLJAu8X854sUGi0kQ+GoIjGC/UMNfFK9zEK3
jQJ6gzlFv3HQks0fMBfarCcZbP3YgPyrwParKN6vUsu1upV/lkpkTRNclBihA10q
sGpRwXszkiLspQEAZJYSc1GsnGczSEYdh1GQNZ4CGBQ8EyODO7XkAQDhsX+hYAYM
Tvep8fdNcP++rTwHUhd6tWYgpNhvMOn1v2WpIQ9Oh3mRn5tFwowyGZziA5ZBQF4G
79OhxEfuV8UAkvnCQHvxEmmFeiLdIgWSBWMqQTdAU+kkKAWY0HwyLFvL+/RmrrAm
UUr3z1aQuZm19qWTnpt/8SlT+PJ9eZ3JutWENx4nc9tw8eGLauGTh42qXAjUNnsl
OrWBZykEFOq5UnYVqK4SYHrT3JsrH5/6lvNRvqTtA7uj+9m1G0hSSzOGaQQOHDwW
KH1rPYeFbTp4UY/2HicsxfIvcdMqUribbCl3dCfKW8nHSWVhIYbVMe9FbgPdgvjS
/TqtXhzpv3+7uDTFU+TFgxRNU5OgkYHkyVd/2EYgp+PeVLDpda6Onwq/5kIjw9El
yTAEkrddpqelCmAnEoP85Uk96a9p626RcWtg9N4rIxwEN78CSDe86gPN3q0qhq50
2ROS9YvagnjDslqHIN5jUyve4BoKzO1vS8KHoDlM5rscB66M75x6DW1KpK0ucZAV
PlPvDk5HreVeonjS3vU7miUfdLT6OYBd7gfyZLeW1KK42uUe6HI5eWZZlWF4dv4E
QYoxJfegfhswqYJa5w9V+jwnMLyFhENfW6s39P1XUxu9cryKtJpQ2/bq2ve1fD/u
g/TGFsAbfSlFXAzin6fzuX3YCxtBXUeoAECJok4zXWhgv7W/4ygEwXqt/0RDBPbn
6I+sdpzZETfErzVY4HvohhVR7tHyAk9MW7iEldU4eYxv2PY7XM0WIV+4UEF7fOyn
XppjAj1vxAJ4h+buJWLorc146PduZYeH3s9eV1aMUlRaHVzFG9qNEH/3tAJHk47D
ylqG4YDo+FjW6O14/p3JlshPqyhcsIn6pJqti4gQOnUHa960axTH6yMecMIWTZEQ
0Rzj0zISwuRdi7n/uXp9rj81USbH35sxN/bk3kMVK9zg+y8HbDLvvmNJThC2eWTa
Jy2eE3AQ/xbRvQCQp3TNBJmmmfQXTAevy8YHduvmx+CrXHt8EcCs86lrNl4m9Lc3
BnN+IJ1A3SB9hBnyU8Zpk7L4hR/G6P+YnghQgRPkebRe6q4pdhSH8fUlH89D04tK
wgg9/P+ok9sE4mEsZ6XYJHz/C2wxqmyA+X7sC2mrZwGz3g1UMnnhOP8rVhDwHezX
IpYj/QP6VUQLSdB5Sfold0BUsbtXx5t6zvG15qKeBzIPoEUCloVKkZdDCi3ZL9Sh
gxRULj61isqY4kVsalRqBCqe7cosx22gazex549ZcddfoK9U7jHnHOw26T/aCNvH
hs9ksD+A8fpnQ4iulgerOD49qtyCm+EQiVpnE9T/X9dKwLwRGTXYW13VQv36D2c3
QEN2V2CziPzLpKaVd3B0TDQZwHLCBdKtS6eOzDh/LKhnAR7XbXRHzKBMaf/uFqKC
MF+ERExm/4uXJbWWhT6o2XHwwadaRXg9FKd6RlgBwEFuPm08qcHPbN62F/08LELz
yk/CZOpztuuox4P7Lo573htwDCRoHGle7tmz29DwqC9pjwzePOYtsm7BftQRZW0n
vP0BeeQS/99INvyggu7cUAFbDkAOR99LCRLKSPgUFPuu7dE6pyHP7e/cX+OomCzF
uyhXPTaCGcSQtkei320bqTPZa/j+HZnW9MRRejNCIFR5/xtJuHh1Rq6gpCrw8c8u
RgDz5CoyMUElxXs+1J61EvXnrEpKg4kXLSWGqYpUCO+qjrNFa5/xvZuGG1B67MMO
DiamaC7tViAmp6sfXLrWpcvDNlLg78ZGu+9ZQbt5pCdejpyS86CfJQL9B5VxO2ua
rkszhedTym38BLlRXakbN2+LgALf7WPX2J4rioa3AGW/rMUxQMqDxi67COGVe70D
S58IBpU4Xk5PyZl+9GJlGK4CgDun3aOn8y3HImeAUL5LDG+ggFf9/jHJahyQLmtb
TmTbpM/K2tb/cGI6PMuzndadhimVcIpi4ZA6yppAdknKomZezQF/TB1WPycjQP/I
vQdMs70eRbmIn9dLp8sjH5qGffeGHLNmj1WB5zHqN6sMuIvHq2erMjlWT00AdQZV
91Ni2iGMN4B7zkRlnFEwuhaOMBnyQ50ntTQUDt1krvvyi0tOJnYWdi1gTI5o21re
4J6DI3IcHuPCEtfYAv9L82guLRSaeQeEI2gt8pYd01mKAKzFlQI0HgYVc/yMHjCt
sq2szsh83LtBvWJ9HMdx+W4muvXWqrE2jfTdRW7p7cMnE4OhJweljPCEmbUaaucI
oge9xlSjFgWAwQlBh6t9dYzlupca6jRgAaqTa+9jpqdwm1q2DlaAX+UwTzBiH/UY
Y+nVKM1GHzfCoVSurO8c86GD8QwuYkrCkU9hzl2TpA2UzoBh3btucRDuMDgf7Nr5
Y5TSBLmB+/cRqSfFr27bl9d67ZHam2/hzXKBCqb2L4M474sK79k5JOekFcfdpQAb
os3DiyN+xpSPPoI634WVKGbVhmDCiMYGoyu0peLbT0rHHKEodmB4bdq8Rd7SS7Xc
0D1o2JVVEZfb3Be7EwzxnYpDsGaKKfONMr9gt265foNJymWpvXxg28cFWHT9q5ei
SLpRuA3eExlebfONZZ8jxOjYDm4qimfklUbm/hFSUUKxqUgtFssjdm6DPPEMOrMp
rU9bE7ZFjmSEmWquh6cvW+qSojSTq4WBrWWXnhe4ZP4dzNzsmGEIsaVZHA07Tnyf
Uv5khpEF4Y2OzF2x+I6aRo+YxTKgyQgg08vPfa9FkUh0x2Fl76Mgtb4CWfN8AdyK
BEI4CuQ2qkHET86S1NnQVpvNMJ4CsxLocsALBgiawIxzTbew81cyNMQhA/C53/RV
wEPN169lTJ8spDYvmivghuxCS+ezvo1El1honl+dMlrf4pEGnUiAn9M0UlovGR+F
wK289SwNnW6iVtVjelQBt77L7W5gO4CFFikevUceEETAK7hxsmO8Xc/865/2Tbc2
hWafm16Qkt4XP4V1/CaIK06Kn3r0JJdRPmIK/nOTHkG5ggQW70FGk6cs/zYhuxvb
0vSrq5VblgZr4FXFxM4k2qiPmyLhNrqOaQn2CB9sY5klvWUPTa80aWMDl4yhk5XK
MFpVtft26MJrUadSQFsuJpedgx+THQxr/UilxFewgg3JEP0TPJhWtu17+1vK3rHK
aSS+pTX3mEt2xWIUcC/8/l3uR5Y4VonF4Jlw//F18PbswbUFAKT/BcCwrnnIQsCb
eNtmlj15HI34+jd+0iT3j0YC6E0dnG5AdgqzkzQawdrhhR9asoxV6JCtbaZbtqSw
rHiqnzZs1HImxn681pnkDgdA0rjZ4lsS1QcPGrsduISkyGcqutu6+e9aTwDGXpGp
ims/ZpEzL52FonWegxiQX43BMF4ARnpZRgZZGdZr8CRxVdMqgOah5NUmsB3AqpFl
uZS6pR5A+wVGDU9vnfbEeVAyMUp8AaQXEN2QAdf43UbDf+YPLof1HzJnWifI2yOR
e0nl6yWAAR4cCuXYjMxQMRHGrSTDMjXqN/a6FmjoYxvj7ux3W0D7yUXaUkHDvAlY
NqpfVUOUh+v5dC6kweix85JDtjOjZK35mIV7PaIfGL9oM4sAytpKmFlQ6NI0Qkvo
YLgOca/P4R1D6qy40hTKA51MtyugR5VP3ZNvtnZHxuzLURNMsC0vyAl6I1j9jBNL
pWLOR18ZZLx6NP6NVoAZFa19byuvJJbIkZ1MqTR0sAnKESpEtz7Gwy/L3g0Ko9NX
WEoMNW8yBK8LEy+79ZN8X4kO7vrQoZWhKQqRgRezHT9tQrcy3+zHltOWZvduiFHu
8QS5QrCQVnN3iCvWCdL6aTzVUjNmhRcEi8pgyej4o/i5khW7Hz4qomkvhnDoFXXj
FiNzoxZAmZPQrDRLdi0CkDpLcuB6H9cO4Sp5eKGucbISs8vDACh0Abay6B/DFMNk
fmeZXfxLmlo6ngaEISW9t54UVq7VfFuGxRbJS2xrJZ5A2iDgQv7HG3kvl8jEvV5j
EAWq8XZaiYSN7QXVdinUbSMthDzgBuEN42GMFIV/+Gsp6VoxRpOdP9XWZeo9sm30
nGVfv/6dw4m1LpxsWgTyzH6z7/XhcnSaZ//r+xLch72Vy+v0wRgiRDd+4407a9jH
Nu9V1rjjkr+7lMwjRplWu/aqx9y8fY2XQWBfO97Ias2Ta/YFUMmtNCr1Mwk1+1Ex
+e3Zcoi7UzsxhGWgQxpvWW1g14XYmh2X284a21ezkQiOO5sTLPGBmhxBjVMPE2hz
fjNw4xsM9UOxQA4osEq8ZS2khjBo2Isv1gjba1NHVmRgUjsdFHEocaTX9F4vCe7Z
4dsdTJ+SpyoOlfspNfjM+0Vcb8UfR9BKY2b6nXiZ5V1MPTt1EQDyDrOciymprHQU
DjxzfoxMnZTwUHzFpbu5fxaIhv1mDe8W1RCCffR8nC+n30Ibw562aGaE0oxjWoQ9
Cyhj3q6WNwWLyDJG+7VMPcHQa7VqEz14eIrDXwS+2x1oWuiqkcreQnTv3U22tuhm
xOjIncPDkx0eU8f+t14Q6qAefUTn8aJkHyXXXSx3kmIWRieEx1HP5Z8wE9ptXllI
Z9J+oo6c0kEnZblxt8tQEKA0NK1bHpM+CJpscyxyYogRycUANcPEagzRTNRu3JEh
oq2Pqx2eRW7op1xcM+s79xutA2INEw1xVU3B2IX6SGVs9vepr1aeUb9kiiGHw7L9
nvNA0uMjfyh5RGsZiXUYw6Tenea/SwwUtGmt5nAqe/IW5WjGo7pyoEEv6DA04ia7
r3sgmfy8bRKVRyC8R1baL3IerdXt65l25846upRN7d0n0ysJBNjUhGZfkNvhjMzP
Vkx8YHnsvnEElunKHO0eLM3cktUbD5Sdi+9V/5/3oY+n7Uop1y3CyGsL5+OeaeFJ
p9/ftt7ITlCZ8D8uHNoE0aBzydvNbbkAd7SdpRjbFopgTN2++FF+WXebRAird19d
caaDJwL5GfYV6Mdtfglu8h1s7I4RsjuG3fHXsZTUVAIb+XYBrVr8UItIPyOpAM7i
DLAQy3K4tcQ3CA3/UuIwwaRLKV/K9Qh9IUOkfpyKf781i2Iw6kLoieSqWA96VVKd
295jSyeike+2bVUvpkhg6fHRDFaF+TR3X4iju0MFxpHu11oxk5l2yR3HMChKdaHj
gl8W6LmCOU/aDSH31DLhgEATV/UownUg4QGoOLqfjUA+jk/wKDwPsk3KxgOr2T46
18QMBhDN3ZIqMVI2Ph3+zIsoDJNaEmPt33o/ILqsb56kut7FTy9LhkCDROZ1PZqp
DjtNjb78IKEnOe0zsl+kG8+8oJcp2cio/TCQQYpKQYXwpDfFxiH/NrJsKlj6LJsW
07XgvnnlnXquPHqITfpEEtdJv5ZVksYYIbpmDLw7Gkj9Hs+tMhk7DL5xmB7o6WiN
qopKwUN8ETjTWaS9xApK+ljUL4z+rkCaprz4dIExEOD72hIebyfghcFnykQDT0wt
YaGN7WPCardTvp6ILcScUSbzgmcum0SOYD2qD6FzC4JHrIbDEU3MsTBTvsXUkmgB
jVMuON0OlTZjhHU08KgZKeiCmBOf8Y1q1WJPClXIX9GI3anZSIDCKBWGrg98BC2/
2keva9qLOUNPGuQG6FQGgVJ3Jx4FlG+cv8Fu+QhGDNux2wmNCTVs1QlYYTjmOl3b
Ez/lFEIQhovchWZsES2RTY57sxvWva6dMO6ZCdZrrcq3D9/Or3rjneWJwk7xn3wS
VJkmM0zplAF/PcJbgFFBVe0sTeKJrc/IifBfCfW80ITJ/tvg09q2c/mqaSiwio7N
cWVvwqNvWge9Dciz6e4YNRsJuQn31GarGWWMdBWdQbdU3IJWFJoEfMXGS99rRPPh
ys8eBqbWSat54k6Kb7mwkPOC9I6tMneMws4cL0G+aWY/t0VoiGoyxOvfpEhsyk+d
eq+CuJy69GkyAFZKdGY/SaXCQYW+ZNNxy6OMmGzO6O0QOioAYC529pTR1LkF8U+0
BS72XjQrdWCI1xAR8ambW7Gli4cwDQwIGU2vMnbwLQsYdJT4k78hWks6pYWTcvI8
y7lnsqUJrOwxP5MIoOYsZ5HHQxcKivFtGRci0oWFmbdDcQRyxL6fw+3M560zx3f7
R6SnZNC3UGT33AMD+2d0FgIRMfPlY6g0CjpcZiQZg0CYNwfrm9fZotvGWV2lm6lK
4zB6xKQS7DqfsPl984s88pzzyUArgxWyHSzeg2lFdp7hIrYYAwxphiO13Wb/6Srg
QXN2R3cGhLisrFhThF4Jy3AUzsu9fn8nqnHBzfY/EtTV1NQNMd3puLLon9PerrtT
kV8bhVQE02cRrYtnBmPQxFSagMnsOxH/Ja4tOcV5Txxj5+r0U/LdHqGENO/0AZmU
lhbyt6c3/IbHEZPdfaIMMkdD/jUMyU3CmJQa0g2lzo/4+BIpVcrQYvqRy+NXa6ag
jbY21kt7NNEckgynzlrYMwNQAkyWKO2XDr6iScOhTLnjiyEpJytZWS2jFHSl47hP
c2DN8Cf1MoypHF494tLlQilo6FpRlHwoSemNo1JHeAYIjo2BUfwGwi7JOwOnWMQU
zGHdad4d78YZWdXLz8kMkHPb8B8/kbC796WUMJn3xR8K0XXZnQruebGqQqnD8p7Q
i1ovcO9OdnbPZ5iAzhFVmorGDGQRgvkrUrGrRQpWaKSVwRboHov1xkzEtRcaLwxh
MQj7fN8xY3j+FjJe2YnjLCvNK8VenVBwLlmBh4RKE+wV1T0qArJbvCwy0DQ/EeD3
/fDybc3mMbNvzCEWshBHvx2XDNigAa74ZE9s0g1MiRF6YzGEikZEXzvJjud+lG/5
7C5ReRjaHQpfO0SuBNqnVHvayYa6ys2i9rdX/j2znh33aEZnU3hKkASCItHT96QL
6h2J+lzzTn1L83dTTufABX30VDSCRBTkuU3NDgutw8FXWE+S+YqD77gyOqA2DhGB
WufeAOmMTG0+TDdJKz3EUPEyxyqwyHzEa4Qs84VwHa+mJqnCNumWQIqjB6jBQDfD
umGHFJeQkvbmhkNUQx8pOkqjc+wtiAD3+lkSH9hvSj0a/++Kmby5hH67KE7Nvspu
7u21vfsOvP2h+ywu3xeT25DV5YJkBK+1RGmDKAhacWzp2x134k5h7OUREa1Zgzy4
314255+qvQyxZAeuqvLIEzpWeNpN/20PWHzv9oTarYTQKRIbcZM6OxpFIdexhxmU
I0G99vrsodNFQAEyGnnxd0jOrz1nDDgBTgv7dh/DWBcC2lXDPcrreORkf/+O0hcH
LE86Pl7w3OyGnjVE62ylODmy7uY8OFRmakiBgs0DUudpTO2lfzxRtnw6F1zL3MJS
5u/1q5xjmEEamwPPoDyktBNExmCG83lY8LV1kbk8FNnET8gl8UK+BEvbTeIP3Bnk
Or4nKI3zjQOgH6ZiGrsLWrqFT1Xpq5uLHLXwDOkoUhYIKYl/IIg5JCbei9ezFanW
DvNAOTU1NdKDyfkZRdfvPePrvHoUmsj503E2sWzT3gZWaYn4zijpIQkrB28IFyrD
s+mx7O8kEdMJQtlP0X3Xlhxkx4YjEtnFe0OQnsnAAO6J9zX+iBMyrTYteWbXpa/V
0H4s2X4Dwm1wxOt4Fkp2K+LqT0aGM5IJ1X+qKNR+kDrwL+abFQA/VKBkWUUmd6HY
S/DFCE/SVCujPTeb6hIEtxnC+0OaVSuBBbe0UrUrZz1wU8veDHppYYWCULm/Ip0k
TvRz4PyJaL8RRMSn3k4e3gHpO57q3WVLHuWYRv7fhIxaHeFe1a61XLHJ8gqMM15/
DTinsMGHazvd46E2XMq6jSCGj2hqH2J1JCWN0kCMg2/2oQag04LO7rh9CZ0V9mz/
yATHl3vsNts2axSFnwwWPQJjYQ0BkCYzile/4IavcyCTVV4yN/fEIWGubfB1mHp3
2VALeW4i/qyi2aw4Ki9ES6Iz7gUXlW6QbMLD9rVfLx/Fh/Aaqzh5SLv9TSXBmxuS
W9dH8hjybt+mbr96rZokDIEfx4wG7TnmsgW8ZbVdcCVwbkj9xXG9YfnS3B3RXq1N
+FWJca2I4ltvWo5xBQJsYagwTDRVm1nVYCfozrIiWXRnbRMdy+mfNtKNURJTSi2M
L7X4op0rmweU7ew3rShBTY2s6Z2DrpCXIG6Fu0TaL8csJ+ICWbn6qggOg9RD1Na+
6b+Q3OX381WOb7Tz5vtjL8sa12lC5erEM8H7cNYAtXvoIuZwD/9Iapb3S8N1xVmf
rYViBDSbrB4vEqY490jGqzRwOlP03LPXc8g2j+BHJr7zPyjYLt1VpMYkchbYJFyl
ZDtMSvzYQO1sTUtT3DXkFFMFgwijJgdR0stnCv4rACNcenAfSVUph9PJrBBs0rgU
ZboEsrtuQjbOE1TyusqBC4TTnYAhe/aNtM6XX7d+jqLDKMPwNg4wjaDM6Tax8kNd
2A4L5iI6IIex8nBCy75oNvNd7WGhrXTCBp4wjff10nmBRfvXIvTUrx/qYMycgADa
CSvPq/UXc/p7d6dueGU6dQPSaA18lw58qcx35rfocjbmBEPum3WRh3WwNarx4BUE
skrIGYzkJoFr9BJBRfWH/HVqNv8+UQGYNm7QcsqxoQoGqkyGLQmnXFW3zy9ZEMCh
7d6EDkTxML7a+T92qZxg9iD4r4pSgerkY7iUqiwcZ5P56mx2VqKpNQM6MijqkW7h
1yrK3NY3YiQeN8l6akHSWYjAKT3sJt7DK7mo9BoURXuyigZ91MJw5f5IkbuCL7WZ
SEq+7qhn92mnsfsWsKzlrrdWeALzxwjCmERIAg2W0WwtKh3cDR4KmKmrQTSVg2XL
SCIqCv6qwpC2TFZ10uIGpFB6UcdZPpY5sU5f3ou4gmOsww4af+fHCRlCvZjtrmjq
PARsaZnMJMPw8f9s25sJNWnCIWV37HcYai5o6GXNsFSHUzFcHj+eVo7+XZwZQvUY
cSOHXP7KIIR0YxHYh/7Y9r2k701l/AXjUULNIJ41MZ0sqNtv2BY/bld67FVlkIEE
pmhvM7e1rdv9gbuNmfPHpCfciPP1z39ejGhe5e0Nbyc+8w2jJSwjIKR0DfRtjguG
y0a9KykH4SiWmwahaQLZdtZExPQQiT12jnY4aM26xMGryU/9DrDMfx9I5dEXGdxF
RLwq51+hkCz3vJNGq0d6g6bs5ZMhaOt7H9AbuyVBnK6YO5zzcmb+lhS6XZiHAFsN
1UMj975H4AZdGjke5RJH2elULJTNTD60lnBm/pPAbx3ASn1SzopPXaVrDJ0PewzQ
7GFXcDVS/vW/hjYQm220GVd8zRKZRnAbhWtp0hRud66Tfa0j5iNvs+ugUvCa5CEz
wY6FJn7A+nekCTEz2O2B99jXZj8wBbJlRrMihIc4lddY8IYZf1Qy8u+zXbcTMq9h
N4gW2NyFhQCN1vAN9Nyn+2OHKzqVvf3r3hf7WC+Oxr5OyADH0agSOgxIrMP2J3rV
MpwlgLv/0JNGNERJ224S2ON53LdHUtrP4zMWoe2AqHzJIVkoYcLKxA7w8h+fgKvr
kFbVLih6PjZ5vTNNycgjFGnu6q9uwRJIXeuOYU3iS4+vCmcOZK6RKhOhaa84qZxL
LYTRhBFxUKWuW2uU0t9KhcPx20mi5EPZ4gRF3f9M6odEHrImtXB0k0mfbzFV4kn9
NFQo2juIhmRoV187abajeAF6KiPbmdNVH0gGM7+l90AwAN3dZnh/HnHOuwyE425k
Vu8zJAd/rxjYxu3UTKX64nzoeXj8KzTiSsKkcaggSVwP2r2tCTx4J5B/Pc9nzyCr
XGIjBeXixZJBy05q5xm4omWvRcHkGGwiYtc1cMMYK2GkreF4yjPdpsppejlPfYi9
OM8iiPfF1q3bV5tjDUzZZvx8+w4AngiK3hLaoGLl1UatG9qSCYIHbg+8HRQpf4hG
NO6iN+sXgnTqsnzVFeJW92uEFWpqfup9jq1gqUWeKwfSzwxMnrfOanaAc0Cx1Xnq
/wXtmLczyqWKMQpHUCxH3zCgub8uVgv5m5t+IRT7brU4Kk/JQ5KCjY+4IQ3+JmDk
qItjC+Lhtau8gTIJCoxCPZxujqjsriUL3dCZph0auHj+clcFjOIEjjli2O7HAsYf
QfJJZT4UTmsZ1BWDDYbWKmCOTyPEFim/pHOox9S2OFCKY6bqvzzCPTRl3mjYPgDq
F9rhKE1r5w3Qm9x5KmHKpCDrLiXYBzps/wV8XOVcHH+LhCWOeOd3nYbetZS0vcIL
Spho49hJABdP0ych4tqpFIi7btEReMWySf25WOUh23LT+XpctG8hMyBP9NYjWMt/
HSnYIubpQ2KWTjWjUBs4kUZSInsz8bonJDzGkBkiFbH0JvMG/Y5DX1/bMAVNdH6D
6vV5+VUrmATEvv5JNWDee6YsHXRHf4JqW5ybdZK2kk6RzQPz1+VyuDdl8A0JNcsL
8Wq6N1toj0je0jk4SXt9EgywplyjlOKImbzGJjHjUxX7bIfHCBtJ/0CYcUVA5BGL
z/gIOE5Awb3SI/SKs4bzK7Km05LLD9VYWlxNd0vPozKEOQo9KkMmHDloVznRVF28
YvFu7uDy3SqhPm4olXR6cioAodZNFJWISq84Y+PJJ2jWi1nX+5Ltg13yGOVWzGut
/XL6S+rZFtAGPlD45il74RJyNqr6Vf6FD1MWSrm2MPmCFiMDU2q/M4MsDS7zDzLK
hdD+rSQZ4VagmzCtv9ulQlz1zAaaE9EoTToEb1Wn54t5N9L+2PvVm6/WhHXG2rc8
2/5ZKhJMLhS0twyu/5w5o8nxQ8dxAOr5b8DNIIEh3lbvmM98SOxEwOgIbhFEDLdU
wro7hHpuYVPu6r2/s8Z+ysAYw2sbKbfWwiz2W8fMmPuo9IOUJIMvr9S9n8o1CdKE
0ANm4zathHN5QGfRJMUWAiH02ETFj2FhNkyb9dg2hBEzN24soAgUVAQ3O4LQPMIp
mEdrQppA/h84019h3m/Fv+aYx7Txpwb3kSnepkhP0BfQnC/4bjjScQ7vbr/PrN++
Yt2WQR8ztkvhOj1+16H3iwAeIYcJcecltMkRl9MZPF3xfMWb7/KkSE72gXgMYO1C
wguZTPaUUsunVBnBTOw9Rl5on/xLja+DHyJIv9CO6LT4R4nmsXSJIpj1deUxuF0z
8w7l2dZCrE/fZIW/bBJCdPJo8TIxco/OHSaj2oWSgJndxRQYLpOVsE4NvR4Y87HB
axG9Sf9kuF67EbP3kOVn99mr8SZM8RiKMejZPUUkCD+frETYKm676eMBudvRV1B/
gfSU3gr8Gu02TQgIUnlvsDn1UrsHn3FEymk2DJ2y3T4ofDApzwJGaKUxoQwTfYBY
6ZkS3s1D9dx3HwzvMPkk535Mwibw3HLP8s+mEPQ6aXnVUC2ogm8y58pqEZpD4Q33
zweoCLdOy/m3KqhRgzYHch0dZZSi2cCFL7/iBRZRLJtlCvTMyLWiHBbq8rcQiHKh
Uy1zEnK/M5ko0YXHf7GgPwvhPw41aDXNtIa8TtIn6GTMWKV2FeEMz060Auzxb8ng
b4WEpejjLG7AZGALDo8Q//uR4f8WAGZVV5Ea5DCPM7kOBFFHeGoRYnBuVXpd+XPZ
kxcq23XxKNWjra1WxZFiqQCQZvVBib7tEHHVL6N5cxCN7KznrZMMOjDS8urY7D3T
klwZm9mqAnhkvS8zJvpW8D1rjEOgIw69YyRUJ1KWMtseLvXjiQF0F1oNOlX5TDc+
fSKVeWETmmTlsRuoXPrgbgMkvyL/dzx0fJWvnHNcqavIBAs/+y8rP/0m55Ad/xql
CiAsiGkfcLeH22sdxYivy7yNvlvhTluE8neJ+R/i7KFuTDg79YjYjv4+nCRKPnUx
D3tlWNpYYOnFnWG0mr5TzLPMH8Db5KnVWiUBKEK5nHl4OvkAsdxnMmI7tHmgjI6o
QbrXMOtGymzvyRCACYlavCwWaJf1k1E9/lEcEiJSMRf7XcZgRi0u1q4R7vIuucxn
HHlFV/xHRWsFV3WutXmp1hgulxvUE8xTKTPs4pkSme5/bzX5khRAC0EvHK88M4XE
hredMQp7EXjRhEWKP65aGINv81iiMSy7TUoJdty6DEXkEciBt8MlH9IZ1vAzwloG
aIcUnzXGKpUAERMuxkYe+z8fOMgiJ3pjlIg2z9t+JpuRtfOABXp38DDRpmaJtY9m
edFWGFBKegvmA/60eYSE9moW38jSIQm8CLZavsyAYaFE0baNhlrChbBNx65e+uZD
+xLgXHg1UhumY74d1ESbvy21P702RFTDOf0sKk6CQRNS8CJ/V6P9F39rO29ZMJEC
lZz24gt1W+UOsC01+h9d//o/1dyEANzrW2M4YCzvukQAqTvPlJKM9X+05NRq1TKZ
l95mf6CjBzqID7qC2Elg/af6ozlF9aURffwih1/720VtscMhxdY6xz2WjRUCIJ3k
tPzTjGuxyPtFnq2NfIkpHHdowURG/y/YDyy9wUthQrnd2BfFeW1Oftt6HyD/g7Th
yFbg+hVkxxgzKDAA5djZLk1IfTvW9ztRecEXO0nn8jc5CR5GZcQVWK29KTQxKWDZ
iO43T82QqYKMKHYyLtGQN2j2BDr5TAfVezxzTHxsRMs5WIbFRS4Mm2OX25uYi5Pn
QkGgvX2zkqJGfsnOH/Q4brbFBzzgk6PxmXp1tArB+72GQEKK+w3Xd0VpvWJTCX1I
nKQSJhDOnyYN6z75SZef1zU2nynhoy6go3qs2sS2M9t9GGH0xrYP3skhooi6gfsB
DVzWhLRxnbE9RIvRs41BHezhKpqr2imUqjoAyAPKa/lh9XpC2PSL2QhsPhY4r1Am
xND07RitLyEI9NQWepHRZP2BvmkQHqowdohAyXPTL9zu63phN1FOtOTUcSrAHVtW
FIL1c3dKPDu/omIBN3NkuXBWQFrCJt3HV2vfQs6XWwIikyr1KSYg4Um2iVt/ro9d
S+zVoFU/wuauRNR+b/9lw76JlaYVMFQbOPkcJeVWnxdRb2vINLCULcPfNN+Z7z3E
svvhVeDhMTuQsRW1mSRSAB9hpsh0upCzlM5IGrHFEjCi/A2hdg4e+Op/ubMbRs//
n7rE63EScxvv1Yba+f+svB/xc082vW6Yor1NPqRGlJgQ664AeyKuEsjdBCA8LuKC
AqG5wREu0aQ9lQRlTetLAWzLjFdmwp6Eu5rnZZK/a57/mYmF71j0FZG0AResfR8z
LAc2xpt8xzbGQ9Dh65NcBrRJWAC222Cx6BD4HfuYdONogBzqU83f/1qhm48DiZmO
FqS3FNAKrp2VudTmxz9HmBSiNzoVlnLnIzXoX1TNf/WsRpykieBIs2ZMzNEpcpBj
67sP8xIMSaDDiMWSCduRmMUfUrGiD9dFE6anrMcVTnfIcmdX05K6YjbgsTumMcxe
9y+Zhf/YNtfVXOjnh/8E5LamSisYQMT8g6uk3+XNNHkqZCAAbksVsAgdWdjBtz9t
ETwFxN3TYBP8nzkULCEtAm/EJjqSOvd1Et3otJ4/K09rY6HWe31uYtZCM4SCl6je
D7Uz6O/MNXH7yDtPh/iaWPVJtyK/Vb1BJ0t+r9/fIPGZGEY1GBPYcjwsZGOXYX69
QRu59GJ7JOcekR9GQ6ww85iX14EuqhHScSMrMxVTYoauORgQ3q6IF1EUpGWTJJeJ
UUHVPQfjvVvB3VLy5rMpv8JraBlkKXdL0Gdbs2LK+bES3QoCGJFEfG8Rc9ikFtLI
CfCiEsd4m9fGDxmUvI7CZk5DrP7sryhW0C7sjzLMUuPADOhK0JZmWsBxb1TPbFIy
tDVZaA12o19eRFKdEMimvUGiYeqTdX+pxn9zQ2T794oUb+8S5I8Fjf2nrLyvxk1D
ASmp5M6rg7llRezf7zCpeWPfoC9MIVpbV0bRezfM+rHma/7exJOX8peRhXld869J
zC3Iyydk7il7eWgTXF15x5p0acL1FMMl3ppRTCROoLfFsaZFtCYRg/+BoqV1nVJJ
iJjhH6278yBCajkSo8eKXm1XJWI56Ts0xV9LxxzQspYp8lj/blqh6xUicrXFeZMp
0njfyK/cE5s6ZrhcRZ91XZ8VbOU/DiFABxKR7GlmzlC3YaD/MtL/B1qxJgGLuRU1
KpXnGE87SJQFUdE0L9+OhnmYC0DdPaezvpcEqNViUyKv/yL1o1d3VvUiB/KVXRRe
gFjIdSWrI8sZRZD/fu8nHxPBIlIgWcyynw9LhPROJyGDH3OS2MxKGH2SuwWU62wn
kxaX1EMRdHHx5U+sKEyWDNJt3/I1xaqDmTtgdJC8wEBjyrlJK+/rP/T/1zSRbwFX
ywIRDJcr+ScTGSyHlqcQo6cYGdhJrEF9+sPpU9xglk0td4CGPfLtG9SiBmQHHOgP
1JE8S2CFOnVV1QQz2KACewqMK8wQlj1Cdbfp4zEeUhYkVqVlJBx7ymrFuc0JBpNn
5KYDqjp7yWiwzBDaciYIitC9h+NRZkXRh0BOlLkherwy9WBs9eKobc3sze+7IPxK
1Ai9F7WvcEBjBh/IwykCmSwggvu1muYG0XE5kIfaylxkvBsxLTUsHyhLZLSZckuy
yXzC7il9cyEV0CcsX885iT9bhsBq4YYaX8sNGHY1uvroVP0JwISQFc0FBkcWvSzB
KKQWpCqTqzmnlyF0PhpSVXVMjaX3ZzB/OI4qVccm9tGHEBJZHMUyn+GSeRlLrq+Q
ZQCv22q1Ad8ugnIMnruHXVmZALy088nXMdoXNQTqXviGPxOUC4SU/y7K5G/ZjJ+F
0rE+EmGrSRI+kFjp5qq/tIfNQJnZYm9/VP0oG5ZsDNWvtq0VTCmkm6ugqpDgbnV5
d4FP4URq5suUd+iXHiQlr+NBH9c7pmjGr7NU+F1QW3TWtX7ErviA9cYTmt4b+FaK
Wu+jMyiN+8giNhAVb5EzHiJJRlFPn5O2rZPmRHr3jDyUbp40UIXDmyyoUTxu8Sij
MDF6MDZZcion4uQr9QO7Q0ZfN5I9GLKv9idRm7ZvxI7/ceSXlRs6yRplScyyENWo
4kuEQpJSJQL4G73zAbu+LsUBej/PqVS4SjNpRyv7aOXyETTmAoiLoOqXUs6TqdWX
a0p+gSYsHHv5TtdrTbj9hBHX4TngZ9fWhIHVn40XK+HwJm1YIGAxK/96H3Jw/BU4
V+a9aQzo18eMkWNWJO+qO39HUh+t4w/HUd8UDgaX8+2oESaAxr+yEMokKitN2WKH
fvKhg/gg/XgWQNAPoaSQZ0yWFBveETQwVUN5z5uS3FtXsqEp9VB8hRQ/Zc3fLgW/
mddqxjryeLEIIIVFvO3i8mQJNNF3RJd8nA7aWyhHEi78nBg+MEnWJ1XMELp6IOS1
UqGFiKryC3FS3ouIMrJHWtAKKIGAKnvX+9gBnPU858z6+VAURg15uP03pQ0NhkRY
RSDsuKOjr5t7fx3JGTXI4hH4LvEMe7XO8A4LywhsKSSAXZ6zFj5bhg9swY/tFKar
oYBu6jkCGd94Y1LQfJmjGyVFRN7XTp6VzWbS0P8+0d6JXrWwVH8flhxqGYYqBmwL
EmSBs8BtQsskHmwljh9tavfzYHCb+vD+BK+ENa6bfDn52tvrNTak7BBHEgFlyWr9
CKu1vDkmJf0+pDN+zdSFzrYGkshcuMkAxFrmiwLJscdcnt/SAPkSSwrhshCLPs3E
1H0PZHoUspH8AxwwW2ZEkY/b1ZpBxFYAZQRfXPmHm7G+O112LUWKCHgXPk04WNc2
Uk2U1B8Qk6NqBT/aSiXjMhAUVXJVBinF/sZzrnf54JdnYWqvpbgl0/rSOsVCipnj
WiiMAsf08cUZpXubyf7mnJG4AOvuLJSvUsMSvD4lVHmCpx0kBb8RpZrarGYOBUay
zh+I0KmAB3XA7JkxkqOU7h3SJ3zA+7h96zRtDVKxDWvpVwmxV7smf+9xR/CcHgyN
qIPWFH/3sPqUOVA9mAsODX2aqpYecG4nbixsnbH7+KVHDdKuQxDxAaAnnkogaY0D
bFaxywaAKoDJsWsy4KOX/eLLY9XLBX8Rxz/vl/5b8GmdGX6fN9tUb+NZmbupwT8B
cVet2TTxRNYKnRTqlKJUjutU5DR2x6Ca0zdxMaBYO56f+rVAm5E2X0m/LXN9T3Cc
aE3Uc0Qj5IhGgUARIgLM9SWH7BywJUV8HbVAMD/jgmDIMqC3igRdOjTGmVEYc3d4
Dv0e/AuzlQFQ8h31qiyP07PIx91OMKcJuF7TK1m4fBdi7Bfx5GsJNuRCB7l62EwF
bFF+OjfLA86PHFVOSBiRlPOxgBIyjlAp8QsSriQDwcwn60W/TByIQjFcrexn5hJ3
9u1U+cd+Stv6cihYTDhzzn4bpn6p3f5N9bFJ1bMKOLxhuP9OZljU2M8X/WdVPj+h
Emme4tTfPFSDlSZHjJIVWpKHObEO94MPDL573Ub4VweyJF0deFCU+KoG0vo2EUEe
uDJJ1ys5F1hLGfgcRbjT0DNZE+RKDz3P4pZa4bvTLc5T0yJ14vQOSZEEeaCvMUSJ
Jx2f8Z2HID0BHdGoanfonUezPL0arnGqqgCLplfhInCEBjPwZaMeKq5RWihU464A
nIwRyMXbC7sF9TdoMfTefOSKmR7zyEAxagqysc2aTB69JOg3c7dypNY5OI6cklSW
a7ScW+vFBdhWj7dRo8LOR9lWHe47YyHpAA9Zzq/4CAC11Xb0ifu8+PEMPc1FRQ5Y
lWbau1VcmKD3Iqp+c4PPFp6M6/SBwY3onoWO44ESvuy67R874GimgxzrHkMH6lWi
L6taMmsyPwv46Sqy3ZVbOVzzdbYLZJwrHlp1r7OZuXjfjsK6cnW5G3PFJyIWess8
jYDK+a2TtWnNgz2MGY+V+EOJq0tOdJoHrfMM1lq5Yp+plyUZKnc4MmC1epPxnRoE
7pAO2lK4L31e0g6XRNLErTkxRQlfJA6qSOsqepzzhPLi3x/wln+4JUAr/IRoKki1
y4vQoCrERgPk8sZEMT5o86P5gE3Agi7aGMsDg98ZWcU/ADpwncHFllgmmETogAF+
vmx2RLOsSXOOghhfYPCNmyYfvwoNEWaxm9Vzs/MnnhB6j7kpo2fPFnjYh4yvEMAv
YA367hNaesyRmq5JRjmLiF++FqSc170D7oE/g3KNSRy8m1Q8BgKJKdFeFZgpa3Db
TFX3JlZgQ+tmvKGYTNt6TTouLKb+MR7gK4o4Vwn/IwG9vzY6s68jR+Bt+yS7J0tE
l8JRsXZpLZZLjIH5kd/k1rSGp+H8+Bx2KNywwTCfxBdmjR/bWWejYcpsrZNWZ4dz
oF6ar1MXAnZe3ColVRDKeODbqv5iof4U2DcxGpSuoCelUSh1x2BBvsoMUfNl0pnT
yG8y2UUXRPvIlGQFHkGL2OYPZ24bTjh5Wg2ZgYzj/uMRSWqnRrnxC/Y2gWIsLJ4l
qDSscnpei1I2uKkh012EhW5ig35OV8d+PnfBpeVc45uEW0arLIyqnFfpJnP9dMyH
k0S9lDXkMS2jpvgpQ0BSlgFniVW6ZkMrHpNBbTUZY1ahsXrdmtMbfB2YEJgtpjBz
1HXF9rGpOvQg690jmCs0cvkTOKUgDYiVTFfI2d6E+oD+4+kEtkBQ99o9vz67+ZQb
BBHSX9F2PBvnE4174Ma2ZFMmtCZRSSo4ecveL6qi0mjdUND7RCAmaMfyVdIuQh/A
ZDIpmixgx+5vIecDl773IQ3iTgw5fuPT2PsSjEJKNuQ=
`pragma protect end_protected
