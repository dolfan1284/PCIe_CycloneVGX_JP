// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OmrnijCDwXcPH9U9X86/UzxPKwM9YcBEmqV0pUstdtFE/iiD2aUDIumhqABtNkLi
aFU9VJD7kgow7e8PKhiyjGtycmnRR/QEvNsUDxirqZHZjkLlX19kqUMuU3dP2rIV
bM59P5KYu3K+NcS2+99OmhxMKnsHeS2LkSv9VYXbWTg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
45Q2YFAXSqHzbaOT1xmcGZsDIwNk9BFN7yhPXWT7lDkFlvF5DuMepUw0HSYJMlZD
cuMOtfiZxa0JcSHI2OzcqZYih80bsRspDjkFVltk5Xyr+YOUPyMTspxHKeLT2j23
kxIt5pa2lZwqjRWpUvVF9Jksnhk/i1mbzTa1iJJHj/pC2Obuwkwfdc2BLrW2ch7c
CpthkyfY+bTSDpBpcxsRUosRSqPtAAJR66eo6IYGCcWuv5XD+ELMwfdPZAE5nMKv
aPhDQqYQYH0AEBLMqqIDag6AzZ2r5yIQz9i/RVaQdtrZ/wAUWTKp+ojmiR8WnYM7
5t6r39QZltSthvuVRSxc/49rPJCF+1ueB7GyzBrF2m5+b3eteETkchgqEpWY2pq8
4SEG0F9U+2TyCxA3YR3oJdBUMsWiRRQLKDkxKPVtfJPHz6IiLyOP2+Lt3ugdWzhw
nOIMgCZg1RBCLAvNHxMXRLzZO/LAoShKS9GmO7RZ/qZuWyylYfyDnYFt1GCtSsMe
Br3wvU5QzHZYM2PYGVuP887Buq+/x0s/weqGRfARG4yV9UAAoiLQBJRh6W8Tnf4h
/eU1uztxm7V5rfmdjDYTo892pMFtfHblSr8KTFMbmjSe0zlSYfIVwEXdFx3gNGBs
vghqdwEEJHOZg28DvYGti3siZV4zLKgLfWHCt/ETOq5C9v6RXHT553x0OeIwXDIX
A3jiedq3MzBsBUuj3xb4wRUgTL/p3l2Geb/TvbFS/1SK5TAoKtnn4mfoELyEYADo
PiKQfHoURYbW5RB7prQnk4VVE0Y3XuZK/Jgrj5JULlK+YKJ2bioy0qQRZ/SwxTV1
YrVL9HthLM+fhJq5SYE5gwhofMB5fXuWpu7l1uow9OugDECVaMiFyUkMCKvzgOHm
lm/Jxe/YWs8rkr/+qnpwcxZRXn6sS9oWdatzA3dALLCzzMLrU3CsKiup70bK0+7N
Z00ygwhnxdl2Xuj+w5DZFEdUm4EeMYnMGmt80KjL+kyD5viqjTClO9huHVHohvRH
xAbLwZXACTrBBBz8wT68hUaOrnS09A8yRZVrV24kaaGr7pPmnK6G3Dq+BdrS1QTB
qMDeOvrqMB9NzGJwH4/jaIQXGdj2QvdpvpWGWaEVxrF+qPvPqYIX/VZUYQhYlUqB
dybaPocVbX9RaNz3CJoBpAvZRZA4t/3BEDEDwGAh3JjoQw9GdPwCg4os/5xSVipB
vyEiDP1f5Z+wr3TCMJQNlL1j8DQICYkyJ4SvtGmnuuOaFVEeXBhsepNZ419/FQmE
K2pFtK/0FTD9x9copmj9RuUUNuK/jyrqCPzuasgLygaftd/SWO1sQAaYjjaVVYsH
V/q37GI5RGTVsTAFp6frsdpYkhD/IOoBa0Svk0Drl9/v29O8sTo0auASGyDL/LLA
sYPSvAz9kjLkFWGCnPJB8b761+kfTOD8p8yL20YbYIM8qyqGSDcBoB/1uuA9fGf1
NTfM79ghhpQrydscSd+bz1C+eBA3/tvJwrdz6xNABgwvZ1DEhAtmTY1g9xsyDeQs
Kpmes5c0CuXFgkl/tuLWagEEh4gRKlE9EC+/5S76msEWFanGRcWMEeApLvC5Owj9
DdsvQW2x/HiDAyq/rrj5SUYgcgRJEo0e7pbXRBg6JIJycM7qsGVDtWXoJP4mmnk+
DholhOce6SD5LbWtmU4uMWuBYOA/C/Zh8tLkNdxxu0HsxOOY6hbRRfFbiQTIOxVq
9Buy1M+wnMvIaAXkHK5AdkTOImZ1aXoI7QTtUdxL4eW/cjpW+oKgIi62GaTS5Gk+
iwKF6TPLVGPcVBa5vIUKLNui+4WL9HZ3I3a2TJxnN6Tl7tNsFW/RV6NJijn8pbQI
/g633Bh70qSnG98yCmJdrxQBu9rlTUwq+4NP40YfnIWPzjC3u+qjV5of2hjd7mgL
mGaqT8h8uCpSSvkEg8T9IMCKom8qbZLWEITTi3nEmDpdoo4+MKMmpLgxb1U7M+jN
qPELc5xnrnhHmtwVns2xx/OZ8CVQdH+xW/WjmjDuqoUwRYRJhE6Pr5pSfCJTrLeY
dvQc9IHGEGhxgJf2bhr9uyQNROWXnhO5RpTXDC5iKbM10iBrj9PbU1W9tdDQOO/G
qvQyXWtBew4bMTD/bbNsYDL1RiBF8LMqE9PZflFFZ8BQnxHMlpaJRxTING1L0o0t
iuQ4BQYo8zM/3hYKSr7RQjMUzlSdv+YUrw+QGaAggRqWz8MgAB06ekO97c0Rhta+
ReXXMH0nJBMVYc8sIObjVkmydcHpz+XpfS72OlNo3EYjfxlbWfJKm6Cs9a/kxAQj
5GlaAnb64t9ZN64LQ/HIT84s8Mn0Makevj/clTJzHzQyrYk/R+LvSob6gMo1+eL+
bEF6t1jUy5ggIBot8qfVzfczsNi3K1T1MB3YnC95FAqzDdOVLNtNJt9PzqyLLBQw
KmVBL0aI41ySTuSn8nOsl7ZDcMzuhxWaY4IBXm1j5/25/UjdOYTaFHxNb6kIZtx+
jrndIq2AbH1Ce3p/JBgnSVVevis5XIzUVAgxC2JAfLvZ0zGA9nT8Mkt5KNj1gkT/
c98d8F42cUP8zJxi2aHC/exHw5PLR9TbFrPS/rERszWRffz7JWPNDo1se2jqqPg/
s6SLYZ0USOFiT0Ti/gHN8EuZqfD+Kom3SJuI4er7aVxWyByHZTedjolQNLaRiG6r
mnpnUiCJ0k6bbuWvqo467+MD/O6m/+iqsPWiH02Fv7dqRgiHl8Agaf1W/igu8+l6
oxz1kAioOdKPK0vGAHHeVoTszvKhWrBdTe3bR3d30bqc+DVdr3/Ua0ufyjnFMReW
DIcmpQpNA7J0N7f+d1Si6++CzPneuBQfBEcY5qUGcvYryNHV45kGwSY2UDIXuU8Y
/tPH6OzTtkVzH2dc+t+Kf9peRkTdY/5qldzgj/ZcFZHd5tYxojGrnvTcx74AOWN0
6BEEKlpG5GX6fht4bkzRAstz8cFN+BXPOnY83TR0EK39Yl4Cj6QZxGx8OAqbsON7
0AZtkMyC9foh9h9oe3b8i7J0jiPDLEQbDtO3Yjt+xNDp8dngCgw1uChXvX00K8jp
oX9+FdvJpNsLXBe7iyjm5V6WPNMqja7U+zYayR5c8p14vCqeHcKtyTTCBVzuO7GG
`pragma protect end_protected
