// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:57 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SaxPgLWC14w3w16kuTBYInMAwR4xOq/m5VM4QYVrXiUx2jJnaldNB1H9Sq+si33P
HZHO2CB7xVuape2npn7caMZEPKFk+GyxDk/QO5i3YjI32U0sBjQRdcNsSpKg+fEw
t0Fgu/HfsO/2zkx/ck1U7IEq1YYQl4ntYbFgmFUTvsg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10960)
UkjCEA7kQRK565J1DwSGCXmh3433qZDlz2ZEgPRBMiTae75lrZuqdAbH5eyloL6V
w/j8IQVLLVYNoLAyxCJov+nozcFIjsV1O2zYPN6Z4sQWK/4NJxDSssWxQV5HqFyQ
m9JjPWvBV5eguNtHfsSwIqGJosGHvDlP3qLtm0nhIgy5SX9n0h7Sgb1+sVMKAPnX
R995mDJHNsjjuXVwI1O0FdtnQ84//HsXZ9uZfa9XhqsudPkE5cj6nrI+BKF7AeFY
H3eSPKwDHCsskG0xpd7d3swessc3EHaKsrfwlZ/lli3IX79xV8L4SBTwdQvwF+bm
+SXQV3/gJEL4xVBfzSXAUmF8DMn5vhfmkDGdEujfGT4KlAFWochz/N2O8mNYSWGp
79EUCbNr74ee7Rs9WGSDZqPs0Wz9vcqT7+bNsT1JU61unwkHbsMHq/ISBsyP5Ths
pH+iDmnDcER/tcTc22GsOUZVv/8mMU7lnS1Cr4kzRtxJLlN8GPbHwAuYPEYoAo59
NwXbG8bfrp1j3jeF7LTSzIsBDYXXVftmz1qr8SSfCymhhk/fVbAKBLyGzRwP65uH
p4ZW7dvJwVSYSQfAj22z3HYNcHqvKl3QlcZKRkwM6zw6I4gtKq8J3PAHY+B0VPHA
zWSxGs+5wrhkurKzgmRymHXqXyH3/BjqcuodbbUYaaLYWmV9gLVgk1lTbOiZMxXq
qD1QQAouMMpi2fGAl7Y3H4vLyF+tN6YuyREpIlZWtZ0Ezzwnu2QqFo7E/JWPImZI
h7B8SF4koOHeOH+y/2Q9p4a4Uv5fDQ5/ubnfaoZDjWKJVil+5ceso9q0Hx7/driM
/ebfUAMlFn5QB+LuDpUIqz4SoIFS/41saypuo+BXkHc+4IU94OR4+Uc6lbHkA7Qw
qNJp26DiM4RANnaXvAjrpSrIn7WqaBTBAmL/SMJnSuN3JkSgWJht5kxks93PHikK
VBFcPkvD8Tg+daHX4hXeQzTaD70QsSqS18Y0CAya/KLF4xBLi3LRcdCvb3uE3O4v
KAywFSAvrkukLI6yEwt+2EzZcSMVyHcPzsm6saV5OH+Pyma1jX/ScJUKZM7x+764
m6FWVbilshGObxQ35w5MC5YW17M1qsbycTb8ahGdxlj5rDskKEBaYfgdiQQyegyx
a5e0DnEg0g541OTJp8w5FavJLJzOHLnUDSuLS/ze4I884tT4nwo1LWgpChzse8bF
zp2zQ1hB/P2zWb7QGvlLwYnsumIJL7LCIOi9UKy1afd4Wq4Jm0A32QWqFxgr/AkH
H1UB9WS+sm2MjfcXcNni4JOEeyHJ/2JvGOAUqqNgcusBKT8waXSRgrbVTiN1YRQC
7PrqnG72sVZOCiIGeNObX7Sk+TGqJ83cEvpyc8fPJpx+wanC2yjuoZ1wQAoJ4oJ8
nNC/wAaryPmbDW7huxQqr44nFUJMwWCm6Mna26vHOF1LmpjzEm0/+4gNKHZtG2b+
SRcVo/CVYxDrCEPd8F9eDfj+soUyRXA+tIxPuKoLialuqNPAYydODDnwRl8xPvbX
HatkRC/ehtQpCgCJvNJU0upKoC2Yl74uBs5qJh2+3DQ39aJMDu1w/ZxyA8yKWXZU
nQUhWjTbGrEcpJg0O33sP4qPrp6R6aEChA/CBHpIIP2juVYEHF/2rWwyBxzTIrAl
jhL+4ZsSBjFkoeBMISELu3xyPYVSYY0KjJLBUwzJWXSt8qwJQPe1kDBKKUnbdXch
Jc7ZprX4DdL+dZ2yNSb9q/mo/wYrrha1n7A5w21UeoTzRBo6L124Ev/TFpTHEC7n
3oDgVWi9OQKNeMRPgDxz7tGYBaTFAvviyHXx459L/o0Q0y2k2h8hb1lL/PFAuACW
N5YcRUI6NhH8QtAr6iIfa+wy6DiE1D8vQLZoBwpeJ+/zHAjkiGnwxprOgV2MX4by
E+ZoYcmW7WwTEAQ7rYtDbeyTJuWJK3ta6a0e5Ns19OBRfiU94OpzpzwB46DFuRnE
2lkbYZpgXile38BvP7XbTAA90+0Vg23XZviy6zmXTGxUZCqoQ56RQy9IFxWWdmMJ
oIRJaDaFTJUcm7+d3FXxEZWXDzfh8scopW+pBredPzGgwmWyWvmyU7353mPWgAAR
gJOre0O8mPF4WYLZ3FD2BQZEnuRAPiNthnnd6L1EMk298C0y/1L+u6Zqg0/K0HgT
RsDdH2tZKUAGmTdG5WmN2Y5UQ1qbLx1L2B/y0aq8UwAodNat1RqNlQ02wxUHsm8r
S7CaABNohfrrBt0GMLLwXapUybfxVA6KRlwqCfluMjDW51em2XuPlvYw8Vz/VO1t
eonH9vslRftDtyakj7HyljElSRBhrmfCl4YfAZSAaWLEVgfqj+MmG1TFq+IIQuoB
KRdBs1HtGkhFLvW0hjtlD1YYyRXoHFGgPYWptK7bH51fWjagzQOYYizOtwgqhsaF
F6EZHD33pHNofQ0TVXzMdOmMWL2xCJkxtBX3bkdTNoHuUnTZgd4HUm1uVGG6YFW2
J5BYj002EyMCHZI2jOhrfdavlVXT2Ovp0xNHvGQJiCK/lURLQc3K3uks1eleNlSr
q35vea6v31+o36NjkUYg5X9NhAIeTNJJjj+hNmDjK3HCvDaMWFlCHwgclh0d6/R3
kOloKCAwet6UnJFkd3FfJRb6w0os1/Al/Szl1HBkEKetH6/KZ4mk8U0+D0QJNycf
WCOaCBLtodGQCBewClmFR+sr2iU8Q+Tpe5EIiyL0VaVrzGeIRogHEOb9fSTP5Dom
Qcbjz/K4rCO3PfLK8M0E7BJmj/fEshVKte1Ouxb0S0OgRKn1NUtiIyIMhYGOda/P
kKKzOL6S4rED9Pc67pW/7TGEpOyM3wpw95lMF/v64M7Yskny/usRPRk6yWwjlVpv
Jr+PdIfuEv3FwfFXamyaIMhPIAZksmth1SNeLJdhjuVs4v8gjYyFJZUyncNImrQU
1IAqu3AwcfLhb3vrhiNYIC6S30F9CU/SmK0uNOCRg2qVgGZLsrkVq544Mpj3Y+eR
A/8YKqOqdSHCHGcdbZqrcSC0A45/cqWVfmdo6pJJz2Dl8Ipz+6/UkHeQB+7v4hEw
icQ24giOJtt2z/gNgl/D/JBAI2LaL3xdOXBPL8KsgQIDW+J3malGl/BeRET4Jk8/
VveQBCvV3XW5aAW+RQy6ip1CIYiXSn9Nlt3hyy4y2rq0rJspSU1+xSko8aCwheYl
KTCIA8K5jIRlGIlQmaOiIPLdMix8uV0jZEFT/94fBZNeFR+O9syg1G2RMKAntCoJ
VuoS6xTf+lR3qkCbb/sP4ThrlwjWZ20/y7i9IceG7QyJIoR7x0RmY0WQYriyUYHf
hd9qSSEq/Y0I9XCoJKJRLqMUlOcb4vUmc3BEqJgzVzHQh+27RYKcDZ8CUR1s0Cxg
k9YbuzqMAXRA9C6DQ2A8SMJ9Cud2XelL8kGhSh2H8X23C9x73HySTj8+YCLTg1A+
BS6KFgPdOnkrRWuGeeBMUB7dapSvVQK/+jO3UCtSZTSVuftQbrzqNpvLFDqpF0On
H/vLlL1g8Lzy9nY7Vexd42bC8ugCupOKg9cNYpgbkVGHm8ohPqdDqdyGheO/OT3B
gzVUo8sDkYYcgi4rhaER4CM+bEaxKCbTbJZR58vYD0dnTayYt+IsBG+leCTLgJ+Z
xZfmsWwraX6Zd7y+HFgTp3B/Cp/7HYanAOTSuOLWwes2MFFYqC0AmwTgmbBAdQE2
RlKqgJsI2QsNIWmr8ooDBLXs60Eh6r1QU+34e4w29iX85OUd6LBKEwJLXVNjbiZA
nBivWpMPhthbN/MJfDPXp66gPZRvPSvUAW/OOXn/Qnqq5/g9EGYgVwzxn0EPr51t
KVPoldejt2ID7XmNByOa/buT9dHaiDLGbg0RgGiAQfaQ4MIHl59jIrQIzbs4gyEY
btYff28C5poLEV9UOZ25CxQAgAf3v5t/I4mwsNUrLBUpAJFsRu6yt8sKnQ0KVQZE
k3X6pT0nXtqeR6UY5s1iEsOTgVzce9Brs145b3So2I6c9cMY8UpEn209UCZxhRUu
dDRj3cg8dtkAq3nsi6U27SZOfF0UJFFP1G/NhvN7azEpuyyUm1JNJz/Owp6AQtlm
E/MuikEvj4ntPtDcr++dxp60CB5XiqCW5zRXl53Cxlpo8nxSUZ/6IxR7zIOBgSB0
lD1CjlL+rk8GUsxHeHozTEsKKpUHksj8SZcAxlpeerqFgCgQVFMK6OB/QO3Ltd/v
CQeYZgWw2sQuhXmFCRQHo+7PPKdkReoFQXChmlmtADemKDXbnQ+qw39WQLMD/nnI
D0E6wcbFVka2cBhi/g64UCji328ejTSYnECkRZKO1N3XR+LzLGwLipGg+fAdEWHr
pydcgXQi02fhe2l0RYWGzrUpj9Y/P7wHpVo7eI/BxTjVZHVjafHUCJPqcPDiysuc
jdWBLXdpV1n3bUIsw/o+yVRzMEnYIFKL0ErrSk2BjNjo61xoj/FOrBzw6EL6u4QH
QqNe0Eh3/qehPNUw9GoK9YUgYi0Xzei0iZwfa63Guwl0XWDR3H4zOAAQ4oztcVTq
mjTJ8O3G8OrV56DORkOgGZ1zy9KR4zivBuMlfE90atCge+4SbLoGXBY2DYlnnPb0
sMv9rACzIDqH1Ru/K+mP6S8GacJ2Ts6C4z0MY+2vV2WVcmeQsIaYLfaX9zk8k11d
w+gyWmbDCafGoVmmXGBHB7v6cTswzz8Fy6XNDkdRkH7DLGM5K7C8vJMnTFDnwj4d
qRUfvVDQrB0kx93EsO8RH0lYajS1GuKrI9d+eFTTMk2cUd86Pz4mCyvlbIZrUMqR
DQToC3ZXZvWoQfXWTLVftjqwLz+PofGWsyJXWOV9eK2RzsJGWcKZl2lll3O3WpWJ
WrUHmerxm1V9NXndqa8jAs6Ih+MRbJbb/dvNp8CBFxbb83g9KmFEKmZJEOo/qAsa
fnpFEbnwWsGSgseVZp6i+MCQm3Sj6X7CJfrReYLmmNhTPJuelUS4Y5PEfG9w4erW
C0YjEbKYBdJNPaiSm9OPq0dYMwjMsaIzZU1YimV5aqfBC/r4z/5wDbigoUtC/Fw8
ytdjUXQ7i9WoCqFhJprVYyzGdneD1KD+TRGSc8c8mvKFCeybQ41SHhE2i7EqkLlM
7qv1mTPolZbSqSJ0ZkkjHW6/FMd8RVAAVTgT5EdpJ6q3XPMB0BV/3p9U6peTbkqr
UQCungzy4GX/OsDtEmFMsP5QpfmZLuP//Od0ws0Z1PFqWvZ0WrxNYn7+ELsuYGlX
rLmJo7ad7yNNTMNvzn3SN+mRLOaJXyHlWr0H7GzT6lOVCBJdoIGqN0TFPJAcnnkY
8r8xvF/imHQMWH+byPHXx9QSz7mB9vjNdSRmVU0KE7x1t092kIadjlUyNX6gwKBH
GLNqG4KSBYRIkNRxBjF3/0cSh98zDfduvPQJv973utF5iq28BA8McwDOz2uLgtxu
E8KdtXCqmnPzjPU4RKMF3md6rtGp0SD2uxEwh/irzAcLZjZE4LWeqglLSmkMTzCR
yGyHgoid+THvVtfY1uWMDI9EE72A9ok7OdCMhXKJefAqpMTL+nj5Fq/AODueJSBY
tLbbfTkCtrzFgxZ9gC72S7evtN1D/5V6c16ZDfTzpqfEThCNN6nxeLugKOdYrS2N
CZmrun1toQnFQs7gYGwb+I5ziVheM/nc3M1vf44mE6lJN2y/cuQBpK0d13SnzdgL
sMY8JJdOl2EiS6KjmCOROlEbTCRlqtgw8VjxhFCgXUbz0USlVEFSs5sBfnU3wikr
9zUJsdUz/1dg3yw2YHv34WVDgIDTF7gbO0vdQivmsxdpevo0cGEOjv7PGQel+0aA
0YFfmstJflaCQXVfLA3E51CnQVfF+AscunQXn4JkrgetYk5Wi3jRWvvMmx+j7kSW
hqAAznQ10RZ2TvQbuo+/39vfJMcoKzB8dEqVn6tqef6M4/XhwiV3hhTmcX68YII5
QTfd2forZ+KXYVWyBxMEmhKBe0Yf+4ys+JjTRERWlCfKhtn+I7sWFUjQ3gTxWHnK
lpgJxqiM4R/hGKliq3eercMWEpcbCqTwKItandv4Cpa6EAw5nSaSB1TZwmJDTnkM
JiVeW1z8lQehUQsmS153HvGP+wo+ZtahAKfSqvS25tg1O0lz8fCITBhZpA0ziaqa
z+u0cvxKOqW2470dcqQziusYJ4QlMhcSKZZMLLMjrW5OCjOuW7//5SD+LRVgrTrI
HlKeV1OFwpz/OpiwYuDRXeZv3NHUsYL478xaVuOYowQshsVkrN4qu/2dtKGwPWHT
kV/7TfexMEfEl2KJYNPuKga2aW90kCYFA8C5XHVBdCnQmuaRe5kiw7X74WLdE7sG
TihZbSRi9zaxdTPoVoF5N6dDVssrJouYRRyfH9sF7/XMWZ/kXU2dlrKzcpUQ4gdY
5CJAy5pnVB3rfeih7w89havBFnyG3A+AvKw36HvdfsyTCXA3cKUNAaJTTfv3F3v9
0+AY953i4VcsxGF3sog131qojHkIqvwVngoTeTrtz2MaBjvk+2ldLtAQAAaxxmNc
pX+Obn2tWHbcDKljpPhXJJ3rd3S1Qv+MXpu+KpqQr/PG+cvkL5C6ThpZC9HWk8fT
QdefVym+LraWoBNvjJ6akNxqxwX43Va2lA4cP1H/rhCnenPq5xP1w/3v/j/1QdDS
OgiMCPtAIV/pNmCbKhkrMSbkAsxsozOHojps0ww0Nn7+NHZElO/LRXgbDwMjU98W
PM91lCckTYg4T4Jtrd97EeC1WFJ/GkLcjuW4rUswXb0Q2fL1ijQecnpXgDEpz1Dj
qNpFytcMnv97fD56iO9Y3bPALw1FPXJ7224JBhpCZVTS1kH4B8Od3wxWX9DwnAaw
TPWUP0jBlv9Yd4fXpCc/+n1dqG0SFZOfod+3Y0/ppfFqxVUPobKjwFRwMKslTq+b
TLSn7N0FFIqv63QcUCfPXmyhz9qsRP57U2rnEKJx6pHLYyuJd2VT/dFnEDu3p6tf
CALGwTCoQw7uJCJ1lACvfQLBAvFAiE2pNKWEgRQBSh4soa5oiDLW/TsFi0ztMO2n
qUgw5jK5n0+77X/oLlmpeFNW+JIje4mQyLu0tLlTrMAcRv7j4JIba2iWQQV6LsPO
W4I4urdZgvZWzq+DKjp3wuwwPTQiPnkk1XHiPaKAK3yeLJ4P5+92oW5RIVk77GfW
ISh+0eLUL1zHI8bM8y1vtQg2HuXaGnAEMiQ15a5CWlOxBZ5Sazm3MKI/wXqyxB8q
29AzuNKPrqA5TCOqZPBG0MT20JDEj0UAsPnrubqR3tUdS6WaxzxHksONZxPodiOa
tAjE1jdcr2gERJuT6nnucuPumxbsg6bppjG5I/rYZm9B80+Jl1Tc42dDBm2yvf3k
AlFcPchDr/5r0G7TbDTtluN24Uf3J7WA06g7Erswx5aQivgsTMx3G9vS3winfwU0
gx//xiNjofuUFQUlITUIUJw4dIRQ/EInTrrVncPXKGPjgsefOGsqa4oeOF2efpFU
e/P1ARm7y18qcX/cwX6ImBmN5uBrn6y6hgfBvRVPpSDLH7W7lSh24h+4ku39lBll
lGY8m+sumo/mrD+mLZG4lWF/6QdUEF4UalPFYeL5lwSVWOGDg3iVS0jUdIz0kLyU
oWSQLZkfiCggyEKYlEnMTPurdUjeK5uomoyKWEYUD2gSy+mFSJnTLVmqgsANDaFS
0jVW+2GdU6Mbn3Am4UcQPoBbiwnJj1aC5jYIi9MXEmGLKuCFxDjuIR77XPLm7KB3
8BMrqRFnK28yqtQh3CtCWepF5AkBMJnIsuMzHSMk6pMNslARiYQjHvmppaqoaGJX
b0Lvz476+VqWLh76uMmWKuat0ViuW+6Y86KpYcXcj61x5ySd+KEfY2hZQfyz+zJw
nvFqxRbisWc1EK3+yOXcaFx2PVoGCKQMV2YsqJv35V+K/sjFPaQs5n6l84e8s4rR
2+1QXe1HDgwRyyy1JOv+RLAOGui7ciWGrAy9v/KVZpxRjgkQ9jMEmD6O86KqmFaW
bN606JBUvsvcK/Edr/4jja3iUHrl0layLKzPLmfvoiwdNECbKzTeLIWUgm3BcOOZ
pw6Pdk0j11Az6aOjc5Fst+xbJjFcU7WQbwUWMa5Vmk2odhNDOIMPqWbpjE/ochEi
ehL/epSEq7GemOPUgC76bfvAzaai7mFd1j7YOJogVK24255lidGmmD+1u6E3tRRS
P64g8RXEHv5oVNfLyFfYz9E7fJcK2eAI21OfyJ92lZuUNSN6+dQwpt4/w9Ya5yKi
bKYlTog5C30j+QJynBUakleZ9YWumo0mDID47f6ygBp340WNrimoI3wo8VB9ck7Z
rzS6+drGWcK4AkT5gjLs+ljueH79vJTM07PgPrweF4mxvHJ3OpFFa333543CxRXC
zG6DhaboeSLblupCBuSHa6HC3X2xm621TWBU9/fAQI3KGTn3QQ32Rk4p413OUi6B
bV3yiquV4jw3/kUn6dYG/4bJIxU51Wpo/QQk/TWWSpAP1kDNhofuapNAfNO4Q3E8
akLl7ghlN+bKPXA3UiZ9v/LN5K9phkHDY2RsavRKoIRmrt0A/lXD95Z/GfsmE6Yh
B9lQP0S7PWIn887Qcdjkm3txQ+/MJYsY85M8oIobonV95D9AtxtMUNDH8T3nRWd4
8uwKwlasV2yJNJCyL8e/0mgyQZeQvETSmgyzbTYC5WYPLKje1fdyZWNgpjkW7LCz
B8zhuFzofV5AUiyh30jWpzPuZnq5ModSm/X8n9yfI369HASK4ACNYzJtkk7uSATR
e8qJykl8F5RI/eauVzLqWl6eiO+Re1rKjOlDG6luMgc/47dtQ5PinonsJoIAxpSU
CreAFWVeHDDvNMh2EoYTJR8xQrsy3w5ybngX9AHDELuBnEyasfx4e+NuZ32i3HNE
eQcTY6IR7GdtpLVyUSCN86/CzghsW9lkp9IeH5B3QkttNqyd+jRDd3hm1OPBoSmK
nRVKJbgawW1iB2Y6KYf1nqaB6Oh2B+ORb6YKR4A+hEgGay2nFJ3x9VcJ8zCxW5y9
VGh28WVBOB0K6l4YgSk/3YHTT4llPhDcPM3AFOWqLWsCOhiEAsouMcZOzZAT/epx
pv4Zl36Ut68qhwFKwNjvc9133Ybt1Enu9tSDX8UBgDzUfR+WUVZbROn2xR38XYPx
NrXUt8ieWKpw8W6s9XFatpTABN0l5rN4JO65+BYveh36kBGf9qnf8haYhz1aLWju
dvOTKEH2AHU+/YUpbmbEJgb8SFN554YhTqc0o5zDsBluAtA74rniYDW8WNBo73uE
Vs/iC5AS5BdCdE17WB6jlprVdnHHcZenKFtwH5bM7JSp7KkaGtU1paxy3+9y5+PX
yCZEaPpVqupHVJG9/y3esvTKYddzS/eDTJ4xODVrmmzXrqud7C0NKtAVU42A0m95
Wwyi7BTQljSrLAiC/VwmQVvu/SCbg0iKah+JYJ1XVem/HQxYMMFyFJ7Sj6velhYB
FW17V0ytorC9x7yZc6aQDKpKz2ppyW5nib29Yj1v/r5afxLomXvkffVRId0aicmi
qc9A3r9qN/gs/aEajj3TLaL2aNrmkfzhob7LegmxmXIF8Ega9/8U6+X36sIGroaa
xx7QsMzbqXXsuONtErFTz99qeEhqXYVJl/aTwB57RmdImz6hC6+7TcXm/HAElx3X
zrFkOlVrhdRf9k9GecflxmcL/exgW7HMnO3zetgCxtev85Cp6YsCcV81Sw+ViOkg
WpQ0YvlGak3d/1DZPsFcQCIx/45wqqOMSGC+OvfbsKG+Jxscx2uOPy14pAXJd0vC
nNGZOqcpqJVtvn3vTzv7wIoOYoBLdwNV2tQITVw5r5590RlQOSlATtDZ7SbVRjPV
Ixz00UGbyhgRTwDpcTkGObDg2A3iORifc4dfchuesZzmCukKVflx3fFQ9MsqWKtN
CV/dXF5Advgj3E4iJ59lsyx9omlWFml9sbhWWOBmk+++pQXJ3ICXoI/dm17Ca4bC
MBnH1/D68FUnit0FfZ4fpZ1JrjnRc3lm+qOVfFr5ERF2NzpOMxLXCGMtfG/aLqxe
g9rhjTz5XDEwhO1gvV7IXrztTGwSpaidLur1vfsHhesvftETTz9+U1o0rkK/VY5I
k6hiQybkYRE06BcD7rQHxlzg4O8PEdcAVWYvJZRT7oQImfwuDmMzYxY8eWuUFTQ/
0pVGjJF4Cvq2RQ9+DJIj4esuV1EEX8tO9QJypzLk4c1x8QvSpHMbwtj9m4MGqnt6
R8Q977t/PEynl17msRDlvHPCLiDbnRz8CH0vOUfOjrBOtwWh3m1qYPOKrlqLaT9P
F2b3F4YR834sdJjUW8RRZWk4BvY5R+gktRUCRTAVOu91NJriD+DX5C4aXJ3JP1vU
8oNAMZUJ2kf/RaOT3t3lyPpU81hNxiQpwWLrRf+rbO4Q4YGgp4iIi5NnF5uxEMSv
xlBHV2cTK452kkO6SCK9WV/zMnrENyS+wiz9bgx5bAUJl0yh7C3iRD60Cg7SSe4G
MXU8yXlPO3llh6K2jquZmuyplF+a/hBxuKwp0p/VRrMuLpOSXAlDF+EMjC6XgDDT
cmw5bWsxbYn6zsGCFPeZQY3CrRNnhi7F0gGm48SvN2WrlrAX0Y59T9JDA64sx+v4
/kaagh8FCa8y1/NFBIe4g2B/FQJCLbz9B1vvCJUdOEoXVqO67e6Mv+0KxC0diRol
hC5PW68Jbwhdt2ubj+jiep2uyTGpqOPmhC5S1mNxMRV5S85zjNDXHmYFOYMfD964
g2LL0ILuClkYImXhQBodc/eDBfq962QDcmLVI/i+arolekirRX2qRp3o/ct7db5x
QkltgSmNHpvy1gGbAfmyQmk3ktsibwFFNnIwd64mYuOdN6emiGhhLR+w4jW1Xalu
icUZHrOqxdIXrimvxzfa1WxI0a9740wRTGO3RoCbq08p1Yk+IfgBy1+XiseOe2mJ
89yXnAJAto19BdxN+u6HyLNA2yLjyd0RZRRUNBr0YM8+P7KhbMxqh1jiD37ihmca
MGY8/xkrC5nlm2/D6Z8kGthl4ZDRwQ64LVOBaXxO3QIidjlH0K4WgNjcdwOPIK2z
9ty49P0YJjYFBYwLwF4EHiRzNrP5GHSUMF3WIyJCGWP9VeaBZuLW15YcYz/phoR5
5A5isoXFQvIhuZj0pkEmHpvCmx0ron91lA/GooMGSzm1jRY+RyBDBk2Hw0xEr1q4
QTHidd5E+Q93VnJTXXbDK6SeX1yUguUVLejwKnU5z3MMUrVWeKAHeR4j32kH24L9
j7FnuIevRHp790jmgKbePnRtf39IsbIYXRH0kjuyRwC8r++Yn6kdZPG0QGYoabyA
/Q8mWL2BQk/5XXmXMKuW6MrXk1zM32TzRV4iWh/DnX8QNoUr88MrZrX3q1UTe+Uv
xGJyyMAYDqEdRYfl84I7dwZ4pu2Q/b6N9nHO0/3d9gqB11XtxZSlPnYVutuR7UgC
7xJpIEEj/UQuITm4/9dBoSq4Q+9+mJSYQ60c4fj3feaLD7seULsCNyCcVyODhJkM
IwmcFRnWs6E+DJDu7tjHCIWcY3Cvk+QApocPFsCYD7dVzVY5r0zqcVqBFpTBdVnJ
h8LNdg3CW5zLWMdq7FQqSOKSBGVUgeyeF/nkmFdlweDUZMF4oyjWdhu+IGWXm9xN
QE4M6/rpxkrjA+wxOms0d58jlRI2UyvRsObJmu22m5SA1q93XWo3vi9H3rqJHeO+
ubmsHfIM0oO3jaRS06yVabhzEsW4UDOImd4jRs7dZvEAssTr950amUKo6lTbilNk
yoLK1XtA85GSBQiXD2lHWwT3uJLnXIL/oaD9ysomBTKH/TFiu0KuiC587JtIqbDI
zpYJ3YbiR+D9TRNILD50Y06/PXzwiYWdeRkMCSxYHEjZOBO3EAP27jaAFK3Lcbgd
Vr8dnUDDukmDiE/oZ0xqOYI0MOhJBEEpfdsKwmsDkWNx2rll2oHojng7LOQRvHsi
zbxUAgV8B43OeOECnck7GxoyyVOWpZiV2TpwExK5OQ4a/zYCncYzAVwTPhipopjo
1MVs1V+P0Wj8M1Y/DEZMpupvVMP60d+QsRR8JMNuT6JquRuKbr60NLSur3mYIh2L
aAAoZHCfcgjCcjmThYAKjycGrH8VdP0PGPjezD8HUQcLPq2WGZSVEF1GMKjYiR82
elmUgEpYtMI2gwqXTOAamBGACtNoERHibo0k6Mv3aGOyU4U+GC1VPvlAd8Il0rK6
0HhAe52FZHV6SjfNjzRmGxYISDN3oMWVA3Skn/d3CN5dSHQKfl+u0WXOC/N89rnd
VEJeaNvSSzMkNAhlRyKkqdzLiSfwzlIprUaerl+AVkK2Pnu21Spbdl7es9NgXXpe
OCKyo1i7dL551uKGRnSGaEw18hifqhv70uGjAt5jLNQwsdubx+c/extHH4+Ic9WB
c6pWA38qUnPBftAHKTNMYMdQGl7I/4Ay27TqIiXpz2Y2Jpht+eziRSHRiBGqvRhx
6JncdYPMELHuFXhzTaUNpwoShbsG/39HkClrFMo+84qlNKi54glyXHSQeYe4kSzj
VPF5aL1rF5fbcruLHpcVljDyzL3+fafAFFJC21nVCJVZry0qItmANIyM7zIiIGEm
yU/nugWG8Ee3eyGApzT1G8TtqkPm4BER3dTpkpS9r5b+ue5upDAmQzjUPUg55Oi8
ixheyyVX08kZUagVtihims7VFSdgZ9vMeisamyHl5cl6UpzX66r8bFwNI7WFEsJ8
rjBekBbD8/7RnMlsnQmXFgAfGUSMyiw6JPCyjmb34kPPAYblKYUD5YWnZsk8E/jN
TOTS8ISwCHw+qv8SSH8TtoHvXds2VPeVSBmSOqYdUiG3IM0in6rR2BQbDbrT1+EC
LTF6K/L1KshmsyCFzPqbq96zqMk/yHhqfzh0JqV5eKCq6Vb5aFhWxuZR1DdQH2Rp
q9i7uf0gKr1x+3wGRxThy+MJmsHnRpVgkyTWr4CuQTxQtCNX7Nepvs1osg51G2OM
/bh+BYtyNU5EaqOX0SYieb7ILuLBTEjBl5FW/U+IYdFNAj7FoMT+kQPyKob4PmpF
WY+SBVIZd06GV1pwX++zhFswO3+i7eQe6fm5TInKZ7vp4eFnWz5weMmCtHQABYNv
o7Z9xbf4Eenu4EFC3jxvH7k1ux24RmGdDF9moLzAbdyeEcd4StmJS3qrTHWhXlnP
p4nAHcEatZuv8oj7z5npCeCkj3iuFHKEE6usTMKo+ppXicOWS9Sos4NIQyDQTsNQ
dO0sz+tm4st7+hqMbzV63O0ohjIW8svbQI24bywVGi75lMMktv/MUI3J6cs70HrT
Zk7b5xbr7doRAlQjQOJOeYIFH2oBDS5CvBQyo4gLmvMgp1/L4lk6EVrKtLTG4H7W
uxuB2O0kl5SOQ8tOqkrMK9uavEFiuhCSzApptBVnJuFMLJJr+Yp4RElT3wbVFNz5
ukIJJQUWz+ss/NsMbCYWB1BKvFuheEw5rP/9leBnnydWeGIeinF/mwJrECnXzxwQ
t2K/Bki5UcJSbbBzA5zLIYNjRZo3rpyOU+mrbkgBekKGdXE6naqZNLhT9wZBCGZe
aogZ9gEKzpQ5b3IE9ubcev0ZjqCLw4v0CiP9dNQuT13MQBCPiyGfN3rfc4wr3CV7
CgdTrahEPpDOmfyWUYp0d5dcGXfzWXuldRKigwPlh3aGEh1kgp/nqoEuQVD0UzpU
Hd+ywtushA/WnjjNgqargXer86CTVAUVtOn4ul8+1x9D/ieuQcipsZbI2U/WEEvv
ASnCM7dc25etVUfkIjSkdFvE+YrNp7QQWsGDvMaxbFjJd49A3dC7OjipJuM9k3k8
QjutoaPBpv4XW4L+374Ze8fdyT2UNedsASS25rS8Bob2qka0OM/BwYWfIAZEi6Mw
4cTPCgf6Lman4cxz6qPzCiAxHfyxsQ/KKyBz5pDEodae12qwLWimOGziKgQh4zeR
Lry+0AlIUjpAnkIgI8i+15kpHVtF+4Ea9HcY2XaJT2V7UutpPfF1wUuTct5bj+e0
AWNo1TZ4nsM1kD3/LpEWyYhIj/jcfPhH+x0UKFGFv3/fRLqFZ/KIbzhpveCLTYIv
V0adSAUPJ+PNz5AvL5UvKKhMK/yBhYQQZPtWwwMTW7ji621Cabm7LSZIYaugx9MC
hdfXTga/stkjR+FyrYOJA2kQvyWaiWx1mCV4Q8Gv7rPKJYpIx7Rzosu+xmCdFuVb
S0nANOa7eXKDEg+TqAN1VBp2+HYxziYghnT8/wINJkNC2VwPqq1/8zV2kSElSatO
A3zIHn1ifhp+TOQC4eHsd7IesWD/Qf9mjJxbOit70OhKgqR6ax4z9JMITyEZfOYD
TXUMhqE5zketrM6SCh00fEODfGzS0zYGQ6IRQ44l1Nn2PK3mSmoltiwi6boN5l/E
VR/TH+UFzQ42/50zdw4a1Vq4X9M0ZOmVYNtWoTHzKcwvDe6aO35ALlLP1VamHgMr
GQOodvlRk3B4lNeYOVbOFh51Dd1WAo7s6eRe2ReD3lVMUsu/y8+bu7YNSEP1rTy0
iOO/Jp2KwlEdxBvUURoyURQfHQZiUoiP0xvc9kJofQAmaTGCODFHeeFK97jRtLCI
Qyxn74GtyK7tgJm366m++w==
`pragma protect end_protected
