// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:59 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CkelcGv7S1QjwfVFJGrepGMvOXx1TgSI5U+/vF6D0QEVjGlxgJ16QYePLqGQ7MPq
vCNpPo1fGLAmyWJzivJVWJTy8qNaYV+p2RgTwOxLurvpW1GVSjavPfJNrQPfRd91
NSu0Il9XazXjHVkTi5UyAq4LdIWWm+lKscWcB4NdZVg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7216)
dZCfmaVJe2vvdJwTz0u61WcYLHO6wd8/78dCXsVjCRK4qxk8tb9WTkxNGqauck0S
jsBQO70J0+jvn41ysHmajRQ80uwLxg2PkSnIO3+lMjqlRJwsoUmWPPdxIcN/VkLt
KT5N591na6gzxW0Yew1F61VN1JIrpD6w/dbMI9EMRL8iqSe0UzcV24IqZCIhMu70
/jfZn1C5G/q02HQ8rK7aQRBxupe2bfGDelVO0+iC0cB781FmxiZ3Whdsgzq25VIj
yJWps1SqYQEq7ePJHdvQ15gBLEOCPth9HAQU7RoJqddr4cK1JQTy3q33kwBJarOD
VvBYMkGdgA5eb3+tuhqXW3iBXylYJ0Udv8UQ2vGljcOe5ZLIcTOu2zWaRoWsT6lj
LaECV/EiOVIpD5OKjCZL6XcGduc71pDug2dC6JshLBEwsUXFIisRt71FHofV1q7E
jCr2k8Px9BtUW1R1RbCwzW1Csl6j11kgUrrmQv0UdazGcXponL0gIUK3xpujTuAE
IZKClwKVLGDd/Wt7Ttgh2iwjqs1z//IwPIBlw/8Ujx4zJh+D3No+KJyC1KoHvnoX
1HEuMtMshgQV39xPVcsh4wehJqmEwszIPWgmAGBN3Z2JLAjHJwpCZHrHFRJ6bPvl
LnRU/Yb4fklNvo8rszEJFE+ayn65QUjvnn+m8rrn9kSvV917oUPZGIFRs6iii62B
RreqCPYK3sZviqWyKP5hnAnYhs5J4is4hSpXuyaUohNE+tC2Bt50M4oIlRSgyKsJ
L3fzrPP+bl3Nqa9LlLoojoUuBRZ+9mDhQ6yjN4zjnnsd0WJ5PyEAsO2HMe/F6mcR
mpw9pf9d//+2zMnurueNUtkeoeRzomoKSHsOyZuZ4/FED07u4gBE8Qy2RQ7fCopl
dMyabBTE1bZwG/geXiqlm7IXLhJTGrC1ZaDJKQZAPYpB26jav7xuUB5799+4G6Yw
7mrkR9iFc7/aP3X1Hl73XcWvIDAIf6Sco0P5wCL5o2JFN/zO0AdFqSYRRGi2UUlk
9Cn8bZ1As+8SwojhY/BTb+AA8ZGbYQOcB59aH98FRQpQWODHKE+YqUPXskqbk/hp
YKL/Jl/TrW/yx7TQrsUIOGmfXQJInSDSe9d+8aCaSV/pGL0rP7UXRQOHPy6U0Ibx
ruF5wD02B57pN5Sfg/3QbIPxbqXZY3wfhmMHJj45/h29wfy6ZoC0/BdtmH3bF7Hr
xjYTUN8P9b8JLNEBISj0TtTRIHl3a8iFNXcCxVTBQtxtCqyAsa7jV2MhEOIdTUCb
jmIJwAShuQFuLfoDZgj15SqdKiTNucknmEShLjdcfSs4bYcny8rWxKqM0fd531TF
dVVQ8rgnWpvmxdlrIOV/Kcctoc4jyf6y5hvirh2awYEDP7f1aHavOzQKZBIZFFRy
Mw5XMIw7VXXfhyIGVgUSwAEn0Uz6c789okqXz36hL6TKRHfi9TyDttAvyAWBVwEb
ONm41/QPAqaLUKTy6wCt4Q4/sk0+kg8hxZmx5h7BBcXGqaAxxE4Y1/nsmPZj9196
no3nYXuRS3e5+JthEw9Cqqc0PwpqLLZ6N8+BRfxvayhXQZuzLY2zcKeNvYWUKIiL
krTk2dZpwm+SJmXrtrjB8WIARiOWSvBXklaGcVsDA4O2fKBL3D9WlIwRngwoxftt
XDO7pUBYdp5tV/zfY0T3Mc09YRzWiwVBFHTA2UjybNN18aw6eelouPzLh3NAWxzu
J7b06csHWYd0nKX8kxuv4/E9LwIsyH34xRhJRQXEDw8tKlWj6WrdNsWPudvEG/hZ
fVKXa9V+oYeZUbWcJsZYSLkj09NVJ74Bn7ORK5JNNMlczJ/wwhGhTRBso91914/M
hxbMIBS2BSnA+bvYtfq+S0Kbsc3OmqI89U0/wexepCy3XsZy60xbJVgTem+qXmsQ
9ZrGpojDsyCHeVlHJmOwrP2rtYWg8FfwBvmti4/wsgWNPMj6mPj9K3NzC4mzQzrl
2hlS4c9IjPTnu8yQzzXMgPXHTErSZstDH5coKnePUc0+dHTTylRpz6xNpvMoiPJt
8j1fRqLIN1WbykdIGn/S/j946axZc9OY2g/YImCBQCt5VnlCI3qTtoFwuJmwI49v
zEbKO+iJnE9cL98lM+aI11veXGeClSzWg6sUGh+KCq0Fm2495njlqSDhwAeTxW6R
ekJEqK6C/T/YnOCC+sXsj3C7B8iwH+SM6Wyg2iVh/71bEQKUBqZk/wFEq/2v0CVN
PNY0NW4/ibIibaOwX4iN7R2DSfaMp9laE9RZv3JcJe1rEcAEAPyUai7BbsIR4a3y
R89CKGH/7SkM0OtRgQLloubZMzcYD9mGooBNvLR4YWbiuPUK7ItuvpU925m/iEEw
+sbHACjS9k0Dw9Z+h+je4BSw3QtLAzpwp03oFoPN9ABe79D3Hc9boiQQFW8XkZRC
kKRfgWNPWFFzk1C50fere9S/2z5FH59G4bzXRtWHC31TYfyie1MM8yh47AG4GqjX
YcD4yCg/XXKZdwFHtnrTrVHFwKlx4F3Jg6dOyIQ3Kfcokm8mK0Ljw7UXnq/OADyM
w7Z0vTGo5SG3sahGInMpgk1BlgQIhaLUMpX7cOY10zcIsZ2S/rFUfRtHRZ0b6yR7
uDSW+SBUBzBTaAIimno8plW4Elf/9ootnP8iBXaMU5ckSB9FuVXyk7ZhahbmsUkp
rXbWvNpX0p3kxEaP4C6jY65JnGjEM4vJhuTqDlHg/Fqk01CRxtbCvW4mzSfobv9H
RyvE71YY5Ei3LTjYivPhtHN6wSzV/QILHqc2vIqrX1M/DvqjAMgA2pzjU7ga0RY3
+vSfaoRlzNlNEn4C4N+0IZgVfySLpODXWJGRDjOIZI4i+WbhXFTbI8DrxMW99egL
gh1y0KNv4ZSE5bCWGn3gN63a9Uv2G2xIdet7CBItTLiVX3qI8hydueGHR0seWiUm
uNO/Gd2FKB1YIRm2BOiG4pEa/sdqIxWVSqtM8K7WDCOS5iy1HKF/rjliOHF5rN73
vcvgcuK5E1kydwQ2DKxQ7C7iomZ17j5LAm8NCjRmj+NQwDIna7Av+2v5QQfjHIQp
GfLIHi24ve5kQ9cf9H9LeSpjyi2dzfKMTyi8SJ24E/bdEL622eQS1s0H8rKr80fg
upK6LOixbMah8XOYpEnXJXYn3KjazP53iJgq4KcPyfmE0CgVSXkToGhJcr7KqrI8
wfkAsx1WlOTYk7UoNvW0lHo/KxyAe9PxN0zw6sCCcnz2gJNZimXoVkXL3la7mWIW
e8gagxeaNWNOQ0Gaei03/dh5aT+DNLGaTkt7igcb5/aOKWrDOrpH2Qi2x2KZTfDV
EWZxYrH0sEpg6+b8nkYumYqeajb+F5x5S+eNxTt8n80n5b9BDUEmUR95GijsHg6o
EQefGZ99Y7X8LRYxDjUis57CowqQ3bhhKdPn7tX1+5El9NlF8zw0ZST+oUv20LVs
SWT9b1Owm2FWTa9To6x+XSTqenuP0DKg8RjIPb0a0aH9Z9vsU7og6/VxMJ5rfieV
g7UlUifZouaPtQ0IzExaR/9bYlAmTLb7T1OQFwK3Fu99pR+Q3x9G2LUUwGG612dA
TN+Hh+a2R1c0HF/W/olyb61I+FU1qAHHRk4W5bDf1y1+4kptFmH7aH3KETTXhN8M
QJ4c+P4AytYjS2yCp2/Q/DBMFw3qIwvYO0ck9FEsEKn8RLiO2oV9LtqEJ706DFVV
bcybXPgPLuV1d9Kf4Mi+4yHj123r6Try6pnZMGMF4cj6Svqs6DfYB0c9YNUV8nR+
QtFLj94lzzGSlzwW7Hw1rZE4FeUAdrl2ZvBabpjw24pwgyJxDoCxuymAYWALVbeb
SNji/FkTWjRFFW8sNAeuuvPu0B0n5PmNuNYYnE42dNEUGL5cP4vkQ9ZbfX4fwn1d
6snAeDnXevGVwbvG625ZkzkV7ch+pIIo0nX+YFnOJf2OqKiN0UndrPGUWSpcYkPU
inKoNHT1Om0z94Nka56i7G5P1QJn6ugjPS9lC9Q2wEG19AvRmx2UJOeY7HzWMsDV
/9NkRikZUQVZKvLdL6K/kE1IDfE5G2mFXNL2eEOb/FuDW30IV7VuThviUv4sa/l+
5ZvMWnXm8O9NGF7Wk1KEveAz5y83ahl3oMkFFxjhh4JJMNe8RnzUX9idocBLpwSd
OcWzSSnaf4sUTepuKIkwvn2Zj+Qvgc+F1sZ9/cANP0/nt/IAdfQkBJ+B44JScg43
5sspJE5knS/nNuV2JAMSYDMG+Pq37lVlxvMNuF2ODVTksB4VZyM+WYHS0sN5N9dJ
g0ZnLxNAOpeSP1ChgDrHcwkI/qgT0gquTcFMLSPgGiecKYb1379DYM3zLbV5lybR
ArbL78vTRPkN99WkpPg7hS1RWsZVF/ynSdaK4cpCugaCoTtdJt/oN+wYy9+cJIQR
gVQdhskXPiW4RifAzBNzuQXTGev18jm0xqM32u6e5s8Mi5Gh+c+m6V3YUd5/vaqy
/QiDI42rO0vR6jIFXu0mkQdcVu4C0GXbAFrjaMe5kAv088Mt24qYRTurxOwrysJp
us0CMKxybroStSrat+zqDKk8S2GEpNU3ysqsBQ/zKWOYuBTbVNQMgLIUPQYQbpR5
drPVdTl/uohaLKce8DptSY8UIMFwrBJk6ADAISBNg/KF5Yp0JWnc0RXNfhDgwWND
qm8RHNXjywXzU45+6oyUlkXjxms85UjsTmIOdbohBztlKg21aS0ZrBYdQx1BKdbz
BSCz069HDQYNKDdZqI8UAVjQDkQ2KZHbrUbCpsjT28aOtgkAmvM9E1pTA4m4Sc+Q
ggNbG08A5vSiVuwLiCDW4wN7Syv9TbBIC67hGkcZ0SmHxirs2GZRy2IYld1JqAAu
Pa2JiqrW3S6HhhgJJeShfaFDCQHz61Bx7Xag4aLgLtL+NvNKbAORBkPrHJWw9Yg2
Lb21rP23AxlTUuyI3pXT3txuGeOrBAmtDxrRqvWip1dutMLg2qSKr/IVce5eIK6k
eNLM13zF2uBA6Om7KzN5dEk05CiymehXkcBED61wJO/Qy0TNMQkSec0rhRfdTdLw
trbSUt/wtjXefojKccc6QT476K6mhYftMcXs2vtvResCkLZJ+HvVihXwk3X84tHy
7qcWwmzJWSfZYZqeg1SlMEKAxSIM7aWDvRnP0dhl7V417PnA+PznaqanZTLDqUD2
DJi7RvQzEUty+ZHCV22hvMqXkaRc1lGfFBnVv8Yyth1GSiWo1kUpQEzIc1l3w9SE
b0Bezh7IobVr/1980aIxAYGoYQzGPGLlZNy7MvGqF9z/uQ8uJIrkXDE43Eq2qiry
J2BPewquVARurIJ9te6zkLzPGh29FJ2wM5+UooqiSo4Lt6LntkFzbTTJmD0OUBQy
YLA69O20d0CtFBQvVv6H9rm+D2lMj6WNy7WS3X5FMYM4MvRca8Xq+SSYUBW8RqWG
ivH1Z4i2+TT9ETTY7GsW6F4JiZZkeSj4X2l5nFetOc+G5JDeswpFhxeu7W2PT+JZ
4jGMwBdlMfPGvPH3BSWQ2J/XI2DgfhFUgMPxDLOOQcPjGYYKZv6queKOgLb98xO6
R3EFUA55TJt+W3EpUkqBvv7/qL7FpWwLHfg8q767famSIwyF+tL1lsxzTu8xl+fE
YFmHwnZ3XM6+ZaPFYasTfXY+BOt0VKaOaOvAvMGdSQj5WJArLhILQjniDjcuXtvf
ES/BzkUwq1qxnVddeN0m8W5YKl8tjBzBEXL0kZWAemE2DOnovrkGb2IV60cDmbhv
jVgYOqroa1hSEsrhUlo6d7Rdo7vZfUZGniUdsFC8+/a9uoPyUPD1WMmGoj/mcpqx
jie4oSMjXD6RWJPUDABFsYmZgaipZ//4YNXvzzU+A1ayW5wHH/0vgY1QREQ4woqM
c1qxOvVRET50owXY0YaipGEbm2/1WtX++WTAWSaWQXI4yDLMHHpA6LxWlSMaRkYt
jNMDttiAMQZm1WJsam9jQCqNb7NZImJlWv6emlA63FbVsw+8N1Aa5FJg8YtDiEyt
PBfYOvmiXdIqC5mK4LpLZjhQNiIMVZICSAnsPoRyAGJuW8ooL+B7hrAk4hIhauvt
NSeVlYG3WM8bDZX3WUdbbXdEFUQHBBJu0dBzlLAIwbP15/9dXoGxVSitOjhO7W+y
KIm3rbS/skGpPu8bAt9IQFMoi6gxuVqkZsoFvQMLGWnwSjbUELsKlenzaJ95lzqU
79TJb7GBoT8Cspgr2Utz/6XE+BmZs1enbEz834Ssn917UDLi+YZckq+iuRvrEs4r
sjpQu1oG1afT67lFewWBaWdvIL7BvKnw81DmQjNrHBUnlbJiGiixS1J4UcGLaBtO
sP4RYgxzr05J4F/23j9V+mi1O+cnvWO+5VVLiE0q2qE7TKxDxn0b9xAE/2/jbbV1
O/WcS890oXzEKzE5jrTFBdm1OQcifiaE23RwdcUcoydxYJf1z84luWWZW8fH1P+n
kUIq7GTpcTILaFK2l4AiZvLFRoZsnARLccJhoiNFUsKcjG9KkfNpC+SsWGJgs+FJ
InQitdCG5K59SkfiLXFCaEtr4UBjTHPmZq7zye89cPS4mkCtxj/5+ph17ld9tbtr
Hq8wZsS9FcJT7J26fwS4xS0Nofu8BxtgZ8eGIRtRx/XaDDH7Ru+z9dd0VLvPSLTR
HhYT4prcSeVC7F+ap8tndVM8ACokhdaIiUJv2LpVO4bStbsBrHWwLaSEq4Js9oeZ
FEfIfiHoGrAQUbvULsIZsQKMejuqvOYk9b3euowWdA09zbqA4SyiHw0GurLcEz8U
KbKzymnURmFCVXt0WaX6//Gh3aH/XAC6y3GoWRrBHsfclQPBcHLib9vHGVZ9cxTz
dkmFysJsA7y+YoCM2Q3bIBdUxPntTEpdntHxv894qoduZ12U2o3tcbunHTjDZUZZ
NzmEpyKwV5iIM7/D4+3r/y3hOpoMHg1UswnlHzghEct2bUhV9i6fTZELh7o901hb
0AvikJ+SjDW9zJTUgAR9Ae3FQTihJpG6MGTr17URZnaOoq0MNFay65fd0fvtQKMh
cl9qsyganAI/zevD56rLbWXh7CIqeq5G7kDuvcr8MJzeZmkY6uOyMHu1j/BdcQVh
+W8fMdgoEkN5mEXV5V6ty7F9LpAcP2Gl+O+4nXOrLSnOqYWYvRXsDJf2otBtPIAz
PJlXHhaDB2pWBMgIuN6Zmt9rH2wScU894JYmn5IoC7W/N9+bMgkYl1ZXFZGm5ZN6
2hOF62+THdipUTqd074NVpGXH5/ZHB57tXiO5UMtnCZseW0OWF53vWnGCGXAA5o/
EZnNamYohGiA4B9OcqE6jdpF/F69k7P2DzCObBsmM54JxjQWotaDbBUfzvf1q3Rw
POdbs2nVYAGSFFoZ0QgHgmfj9I8al5CW4vB9+8m+oZtvLV5z6aawbNQLNvzwZ1Sm
sm3irWkA2UUmKZ5eh+64IRvqx0lbaeM1SzFfDs40uaQsxTyKZ+kRkGd399H1d1fJ
ijrxnhMS2XNojfZnyP30xzCCvAvPmLjTUBtrNIkVfPkUCn2r4MjVRs5RRV+elmVw
EoBPExHj9WcyL8TSzhT5871+T28eycRrj3zmCjrc7RtDbzlAvRBniYJnyPOCSX/I
yiUdgAWM6CXrfk52fl1ojBNPMOqUewATe+5aNd4rcwdW+iYKoOsfw67NjiazpVAU
fOX6KXMrFGjXmqfyDIonrmII8pbK+CoJPGtf6Bp5d8WFmwXfCRJmQPqucbA/oC/U
uuxuBdM8KiZ1B8BD6KmmpifGiKnPL1rXc00xrkUJhVp2bkU5YtS3IPipig/XuVnR
2//SL0hZtWRGmbJ6gK5Fxo6YrQe6JsxMB6wKqOGyUDkwlLmAqujOQONs6qdpAldM
SEv8t9GKSxS/IcntjQyHxMRrnw6EHyKc9kfnWsABq01sGMtX4QFDsUO67IxSBV7r
Zq11qzGzaUurfsM2tG1755hZ0M2KxllN8BUrpMIYJhqw59bUKaAdjlvStXE6gfJK
W6SUeFQUWeDu70W4UlbMU5D/IqlvqEol6GxURSH/JkGDODBP1t4z56UlYiV0AX4M
vnRivGg6JU13r+h+hhkllOyqE9tMcyn+9W+g8ow3z0eBvozzJv27ymtmu+sx6k44
EGaQQBLRIMpr+yRkjavkFhMjGk/4cYzxlRlDKIkxVoh5mgFlLOWoVvOV/up7QsnA
SV+Ps3SjxZxjJw6uS1KeWomTXx8LwobVqFipAs3YzTKBB6QYkGmU8Sq854q7HUfD
s6prRUDM8p1z+1QPUjQNB6/V/cfV8qp8yTLYpsFKnhd/Lzw9SWBUPROF8k1JVKBq
0z2M77I0wfecbE+O5wIwc/oK3W7RK+dtbM9YpYFunMVPbf3oHUl3RT4ixShw7txC
/+3uFqSE4JJPHnNBw1IJizeM/CpYqu1FePHcBB4wKq4rEyH2Yjl6fKpM/RhqfEgG
nuTBtXaRFru/cr5BdckvoKow/IfONtJw83CF6KxV9qHuO+CGis+kDdIKgk37tFnM
LNKto0H/BTHwJOE5TC88AEaF4rvqfRl+QZv3yYjomdNJZ3FQ3M+GRM0XgGQTUQst
RJP6+SmmiOH14P/AzwrktFV8feqkZp7uSY/6B6WwRjaKW4103jfVmbs11x+EwtCR
XJFoAynhWr3TuV/NRILSh4FIDIEVEOvxz8SmniuUZuADgtQUvzjPp2Sugd6ZRAzA
yiCmc38DZOgWwfDrpHIhGCRtURVu79u/nfzV1AyRUAq1Sj2ID2hE4wBLgeJ5wdbV
R9K15zjHZ6bVVjW6JJ07Hhu8WYHD7T2vRhZmp/M2PXMxbluGqHQbjl/Rzo1VNyYX
/tgBAgp93TdRVvvA+qryCJpSrCwew6xNny9h+X5IuzFY/38yHJTTcm7SbUty1HU4
Bq3dzP2JpHY8ar4bqXfeeD/+6UNr+mv0RmD3cjXpSnEvWsuxmZoMpPa8ZkQZ140u
VOBuQycL6DpvDpFi44OuSskx6eTNUQye0H+xUlrQ+LsWl1FQUyThtRe/uEfxIELi
nY5M4514f+UL+YdzKkqCZx3CIr7Pb5ruOzNL6h61DOve0BtsjyglX1NnyhwLP8MX
NDIDdS48cN1WLaVG5XFTo+cRwRPUch1sD1OfZsewYTcf/Ln/JJNP2KexBlaYiH0W
/ZsgdjUOQteJFAjjIAbaF3tgD3Qi14jcI+TZ1I41hQr23XD3QpH8b2i25H04CJSJ
mgnUlSCt3sZxONUrmoVwCWI7I3dfX/wdhfn/7d7Zw5yXGNcHVNbVQEgYSQs2srFI
Zr9S2h0avkBBDtgNMbzZNqWJNNUoh9EjDK5gLqVsRHoyYqMnq3/aEj35Ze1wUnx1
bfD3xTk4JJEmwemQ/e1j96qcXBAHKYA14aXeK9jNUlnrMScbu8nA5DFckMAfnQhO
v9GTVZ+gX1cyFv700apibthjcoJDWdqnPj/7Mz8WHfyChiw2PPoOO/IGX7fsXObN
LpjPKmIkzHQH+VJO3jwf6n3qq3NJzirC1DSPEB8ihvlIqJFfZPu13LFGaC9P4zW3
VT6+Yzq0KDGxcb2q+GtJfzy49JOmsONgPoYVzRr31SytquTsByYFUIlVqR8bndom
QMY7GqIdNuAig6ddKx17vw==
`pragma protect end_protected
