// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:01 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iYgHUi+4RbdK5wh7ZNCQ5qReNuBoFqcTxdpHSSyo7RRwVoIn0Ed5+NAKgygQFZ6q
DYfiDoklgXF+1A5Bf/+ElhW74XZAB71c++cNWqn1JmtyhYVlgeCQo29T9TnmGyWm
pRh7LIossi6ZB1QfcIojXuhKGAjnFlMNDuu/fKSCQFs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3600)
fumFn17kXAtk0YtlhQV106Msj4O8xXQSi9jB1K9EOEBC5RB+8f7+pHmGMr+Ov0iG
05iRdJgV9VUr5iW9YUMjN8uMFojQJKwcLX01IeFJFQ2yZkDKRDSAnf4a9Awozlx1
tv+5JrGTA1F5o1Op3lz+kWvIGFEuyec9GAMaeW+BBMb776qRLQzcZG78rjQc5JDb
sEyMiywGqCqhYD9QSrehpQJjGZK2LOtxNjb0Dv+3xHN+laBVmFbDMZNr1brmdmBB
XhQly+NORbAu3SiVv10NVh5G2WuA0vmlVcDTIn83NqGAsm0JEJ2+e2y0AbyCXU63
Ec2Sfm4PShVBD3mK8y2dIEL1nGF/GCOmei++ixJnDrUSzdopLzf0xkCxx0BgiaU8
TpS8jMuBwxXeg0jG0cU36Cw9Uin6Bpfu6T2i0OmmcIsFGeRS8IMhQ0547Mvby72E
ZSWseaSEGbeRyuH01niYsUCAoLDUA2IXRC+VHMR6DlKK14bTMUbqjsLCBGTCprlJ
4QPmti+xqURjLVyoiyWCAzfR3lKU0QQzHpJ/bUU4lM7eM7oNUChcOHclXN9tLKH2
587hprIGwTSzCjGJU7FcAdxoiHPY+5lanwmjV5zq88srrJp2nwQimyzUv2FlP6jc
NAfYt5iw3UCqYOludBOkRNLFyp/Pna2YDpqHpn2E9ofNku+rZPIByFZ+SptWhOVH
8FDf7N4HGc3nlDY8sybFYKaim9ZN8HW6ZPLECRssFi7MNm7uZveWbPOV5OgFP4A3
do1eVs/W5iG3fSXO7/GIu58XrhLW6PgZuPX7mmIGqRKID5YepcnnCyKCOT1VcqyM
Fk+q1KGzj5VZulBdy1UJZ83KDsBzJkkiBavkUODIpwzgxYR6o3ZhYwpBCV45F99u
mOFROXxlZR+TWvmldjkmdJTf1Axnorr+f9Xvz4QA9z9x5DS9zHnT28TnORY4uuhv
ZNrHntpsiGAFIMDrzW2xW3B0sfHNLbMT/PmEGza3u9H1rnwjcjseXehuL69MaTGJ
E0915XJ/oVZEf6pvGdemDAlH/D3FLesvQnLvKt1122C63UrQP8hDNmA0L9e/7rao
Kb+ieOog3vUXBzQb5DXv2pqN7KY9nsu6MeYrlpxGflW8o2EbiD1GkKX+bwTo9Bdb
IfJSNP7XkNMy2XJy/nuu0xbtAg+ezDrCFWaF/ZV/Ov9/AHZKwLBAHcZyaBQOuRnQ
b8ukAZU9zgQ28nFahBbsiI+EiJBfFOXQV/7QLnut+MzdkLw5lAEIEsWkzJWzMf43
rRr3VCOZY/iygDosIbVichRd2nVjMB9TfJ990hUkgpvFE3bNsAMGweZM12rvSZPY
UgAMutdiAyc86hVMqxWk5n+jMPxlaVlmHQ2yrAGGXLRy9vmmJXEj3ExGv4pWaKUy
mXgp3hxBLW+zK2xjhO5Nn6G/ZijCjJE4J8P1yw+BKws6ErNPUZTYg+jlUxMxY/eB
82IzvyS9hq9WJfC5Zye6w5CSLX8Kr2/VxqRKe5/HijHGx/LKmZOp98ds5o/XyHiW
3csz5KCiB+yFDdW6xB/hr8Mz/Z6P0OLqjzekJoqP5bQhZkNe22KZMTAAS2DaYriV
2EQjjcLTs5WRMnHjN7mWsyAj0rhkoewL4ZaqphY1Wkz8EcS30WLeQaQ+xJzr0+LW
8fnZA5TAzGkj3xzvkKFcywzyF0kFuVOR2fgUQhfJgQp4OBise/MlBOp/i0psH6Hj
/2NWfq3rYXl6XxImv5NOYNEgFBHDHFl/9ukTT7h0UAqKtJPXm19w1lJgoWK8BvfA
QHg+5Tkgy8q9kwn2XG8ImAjtaKion6C3YyS/5tX9dizQfTJyniAZZCN7DvvaRNeD
ZDoSqboYXJPxeqELVty659uQtOiDuegKlouBNGpj2nN9wSxu32t4rYjtFv3k6Oew
VIIHeEiYR7HmC3r9bEwAe5idlrM97yKVilw6Mn0Bu+R/OJGR3WOaKFMVVIsD7Zlf
TlMQ+KlGjsaRUO40mdLFmegzYhoWrO4hr1nmMsGP6i0aLtc2rT3/vBS4bYqxBcOD
C9cKRVflhyGiH+JK/9zXewqyDgkYBWylBbY2n4w0E+IPBaNLrHhXqB2z7JGZ62kZ
VY4OnP5s9LVvljsigM+4sarwOYU0rPdCK82/YtZWZem2qzIYiUcsJLF0YRvKEqCY
8oPl9wQE5SdNP4O/Aw94cQU+ROrnzNCvhoDpTQVI1ehNJxheDRqGth4oORIg0Y5i
BWjmul0xm2J3G84zgywhKKLFTVk3WCYyPhU6lM1IrGiipnnzVZrlDlhx+tpZvken
vHOM9+raKPURnLXLPJiWyLr6cy2XigAB5k8UF7dyIF5bcf7ciiMIUGBj/jXvWf8k
7iPsMGYbZUAsdXIEGQ8ArFgQLh0vVnmOBmzqaPIpcPiyZC3ZtlqTDOOYChqSED9g
40prBKKbSYskGRjrciyIzSr11nQjxKAd9PgxiJ5wmySkMbbmCgVGf6tZekzr2Xw0
GSkCt9vXxIYVQd/ui5c7JpXNZ2QHasjk5fQm79Yx40u/4U7SG/aBmO2gIqv/77X5
NYOOaOHQAn8LBpwidVXeGAY7pEFQB3vfOdxno9jySvwLkLTOnO2MS44iOs2XdxZD
5XJjw2h/sXvBhyQYAp8LpayiuRtdy8L2A6PiGjlAtBLWae1azCJROO5Q94+Q99+j
EVMzxz1gomssEIeOymXeZycH1yClT2tFEQpCcC1Rz2XVhP3NTmG5iQYdszzKeLd4
1mrSIYhqWQeMHywXG4KN5k5kc4MSE64+YlDtBWJZTIc4oBCky+msr9Aav1vMxpSg
d/UqxDTwVQA6wt+k511xd1iv/EtbHqPzjUfONGWQ4Z5qgS7vj3F3ORNy+fiXtA3E
h+JEcqUx9LKxhoYB9heyUKNuNIdMr5YtRF/fSRfAfkMFKAEXoiyezcqLYGwX7JSN
Dg9AGSE2P0oI4sZ9BQ1fYb8sfHvJ/E61XosQPyGtw9If0uAdYES1pSB3pgepPO58
CBgwNMI+0pP7MLOLKWIlmVF4TS1dRwP1h/Cgb51M+WARagf04+36aBcUySEUjxva
bg9grVm6v9V2DvwWuCNVddvQ+0Sr16zI8mbIxwM35UqMpkmH5DQOK+H6PlcecSK3
Qvio6ZD94A4K9+IHAzsQin4OhcWfZmXdIZY72nadKgVAxzMah693xcOJ2Y4XTqIE
4pIsEdt8zC7kJyFOi2mmAt6s+QSrcgzON3dIYYgFkCKkajhip6tc7woQBre1paD1
HEpADfJCGc5aiB68+TocDlxGH+dLHKGyzIOetDfAB6knyC5dkFv1J6R7Ff0fKIVH
LYN2mRSbptqXYD47vddQeqCo/HtwxK2GVbLwgYPil7jJ/3cZvGi+v2WKYp5xDW9w
quFPX3PFDZOOrPXamAYO7eQRWRGSAPWfENXQ6SIvpc66Qvb9wkQEpKpnYd5+Zjpe
ltwWy+H4+hABq8W+sk65+5MgevmoJTuG6Ni1CjCqTd/IBYW4YXm21Ez6IyuLwLUQ
XC7WUFhrPILg7jc1gvk2rBwYjRJltGuxhf0Zep4t9sIOHsSqJEKSwg5K/qLX4D9q
OkUzZDf9qlxh7s22SWX1ZeJgxXz68omddi9VToxhUkOtz5jPyP5KE8EB9Hko/yp5
m7jXYpTRMpkrLE+JbCyG744raOFPlekVK0PWPcNPtWLz3WkZma2PWu0O91uUT28o
yDqg6RzDc7RmLj3Wse+N7/EzM0DEoF1+WDAMNSnwGvWiHII4iT/bPEPAez/Emr9T
E6jyZk6i1X2448mieJfJBKBpzdpWmDe6iTd4R62ATQxK2sJ5xZHm5Fg0gfZvwX06
toSk1GBReA20wqYV5gv2/kURc/MLyTtngSL+frT7+XagTnhXN6tfAcGxI2Csf6yq
UaW1CJPG3oQiI+PX0VyZGsMVGAtekRl728THZq7dt0S+yVimIheiijRtJDoDjf9D
oEP9k9lyTEAows1+ZBJxIuE0i9QsreXni6E61UW3MkXr5LxT9s8oUXh9tHQvCcPi
sOKLx4hpCOFOEWlaOHSBENzW5+F54mq7N4nORw2ocBrZ9hIJqNiZ2cHeQuCVnyvy
HMAMbO4OEHXCONq5tlw0gVDq+Ipz0PKYLiW6pSbonBgdq4Pv7AMD7Isu9D1f9b2X
vJnC4lVPRmMu8FORhWMLmkEoAlLAWBbAtcSm2TGeyTyEPnlU0q0yY/UIHeO3H1YI
MOrLXMSwgXTWbOFESqgq8oN+eF9FXF0DVhYvxmb9AkMxPMYKFnzA6GP2pPfZzelw
5hEXJoQOKZrXs3oZSyDfDn/pM2/MIBhmzJGq7noc4LWkNqeKA2g3D5KzpQPMd1yY
AZbl0jinGant+UFAvqQI5gEP/PiSyUkAlKL/YZfuCRe2klqhsJ3Q6XLEqcDFQydk
I9DTeVrgbvSG9hWqad3Zn+lEp3aspydXoMVJrHK7ncPmALN5DePfnBIGlFAhIk0Q
zvReKrpuncKCjGRpnUpkQf/eUrv2EoB9r6vMRhuwbjtdByuynatTzi4xH4XAtdmi
0yWMZiNaFambTPqPze+CgIruzeRPp+rcIf9/j3c78EJB5V8ZwFe0a09kpKTTud8b
3Ao+VuD5Ty7/XjMjHdwvCapEAtL0lm4F0q7JinsroNUGMN5/RtRNm84NZpUoLV1E
1JSwcHwGQaW9Ftb2iavy+Ea5OygXDuYJwJPcYjRQ6UJCvHILrXshkNYDCGidZvpc
50rzfzkLgVXp0J1NWlAR17ThXeTAWwJosR1RKYyT8hHC4PS3gTxnhvNuEFMAGOHI
`pragma protect end_protected
