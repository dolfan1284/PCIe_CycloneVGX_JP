// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:59 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b8+fR+6QyCbBLb9yKpzO3JqAMwtxiQ19SBTiVwPeB6OTvX1aZyHScUkyFCU86f4I
LDIf+axjwqjFVOCSyUycsZKi3stVBSLak26vYxhkDEYNl39mI3dupkdWc9dtZfSG
k5IWwTMUZzjAr14MtTSi/oqE/1lDIExnfpCzXf+FeRo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
oQH2WYcttUjD0pK3IEvCQ04A82p/CXQNK3AxwmKjTWSbWmjXjxTV9n3JQ6zhSKbG
RhPFZXtxXbUuLoSK+36kzl+cjW6VXdKQbDJRTpydz4T+UDK6x+EMoH2lDs/Wo6tf
v3kDryk5fXMp/kO+x3MGHSxwrXMyPHw08VVaKuH/PTS95GwSxzDggM4ljss6+3Pz
zK8Che3e+M7/G+BcOo4KbKq9LOYcowczc0+kSox5oL8u3ok+XMESJn8OzjzeutzX
xVA/gXxT/DB45/V7UYPNKdOTX4MrL8ZRSUdI/lEPtdXNxBfN/tC00lv1McTOlWMT
6mRxQMvv3kpZxo+CJ4sRsZSfNPls8d9YQlccQ6O1BIZA5EcXZ9rg3xkHfLjF9OPg
pDCBc2p1gvONIwKVk3kCrm4qGZWR5v51Y/v/I+b82kJtPjYclNMAg6eveVBj818V
abBqMXmKeiQRNFUYcrafuc5YP42Il0kf9TeXFG2L7o42xh6LRuKHEUSzsQQotYPr
+EfQdFASw0oEpGHHczwh/zqOFWXOCV7vr5fKAe57ME4shzp2HZDGGHbl7y/a9fUg
lhixDichV21wo4Z/i8Iq08sgD/rP8sFfDmOYNy+Qrs9O9e4BGXREPBqyW5S5+87D
Lbc7QsiJpmI5qSMgTgRvWMlX3IPrlRxpk9h0wqFQjZtb1LFKmQzvaW97905W+rIM
ZY/qYsVitFTzmStDUuUn4GOdcitZS5HTMAs3WR2PcxpTv1KTwnAkOkIdv9Uwy5Xk
e12RZj14z4hrjP40+j2IFimqyK9+PaeXoSK1nRblbP2Ywv6L+Bm4dJIbWvpte4tH
ov58J0k82fdz/K/uclGQRrpRREMI9MUXI/D+uRulk1YlUy5Ww3Es7fTVchQQjZXG
tXuUWhIzJhpcjqB2lTXAX8s9+kpYHDItvgc0s+xtS4vb1966BCKx800LZIB/xa1P
FHkdqnkrdGjMLXY7CjKb3+QM7cD9vH7qGKnXIoqBrlm/TQ4ayOEWX5jIvAfQPnm8
bsltgDQhdxG7XIHxd4ocHnQercEZlygN5B+9ZMrzHOmIb7qNQvzVUnSQV27IOh7t
kbBgqS5cZxU39UolG/TvMuXnkwagDkO1Hxbrc62T1dJwml8VthdzTSEj6p5FZRWy
yDiIM4/m/zOnQ2W7lqGg0Vs8Ahfns4MYBRbWxXvfvPTt2PVDT9koVEc0+D4MsyH1
KHru4XK0RcFpGrJGNtKlBToadJRO4/DIm9CeN4wdrmt9gFLYVetoFm1YZn24eDxs
4yFsHvNvMoJb/zi4Oq6fxXpxjMdZ4Y51ZwoPAnxUlCh2MQoy75aJWVwCRvxvQPry
89JpcWBqYlV8ccM71mLOkeNSSyFUFZaoLEE/klYq8nF8AJH5BxS4JAlAAg+Ebj3Z
7dgXdR4eJ0M52Ezxxp6NGheV8hiu8if0Bvtzo3kgvwYJrqOedKsJOH0wKsqFvCVC
w1oIusipVCQOGVtgGj63iu/ER2h54IBdJDHLrdzAXiR0NJALQZ6rWYaOwNm8a5+z
AnMa2k+JjuZX2xbNf8H6KJniTxkmgkws2U3iDpsp73yykhdkP3718vQtwFPoKOEy
d0bghRJJWoyLEFLYoAodduWFxuDr81v1F7mkOrXZKQuN7A4Eu4fdQMV0YmbZAPtf
Kz2TAzZ5NwxWJ77Rd3SLM5sjnCIlnSaw5CtB2ZgK+jar+NMud402aAjUxZF3LAVe
2xpIuMKSWIqP/NrdO3XWb6ZrRGLak4RaJW73FDRCyuFbVT1SoQYSL7X8KAe+G1iU
oBeIC0E84FNAPjjF49qnZ/qXaipndY1XRSXphyBFcJH3WkhFIj2+PTwlNTtnMAJT
aNViwmhKHwhDCWrbeCgZV5BEdWOftI2bTl1U1cTv7+hcZw8bh1Rx90D/vLxZqgsE
yG1Z6mB7xWSlsqKcnzG/3ufJsNKDXWyH/ExDdWcdkkCCy0ROsE7wUn1hkHkx+CZS
w/sUgN5NIs4CJwvY/tQLGYtLKxsC/WFEKb1kb5wu5E80djpPF514VncoetH68NzA
dm/u8GRP2qy7g/oiTujD4BdISKN1K/gebu1WrenGHmp++fMGL0nH8wrO/FGRJ7oA
7rxxrgjwmrUWY31fhv8alnyhq+8+L+srzTM8O248ZilhOJjHCWe432zlTO6dgs14
PoOCCsU1sfusrbf8suuQbZ0ks5na5I9Ia+L2RFro1iTV8J02AvJKP61AwMtXz7rn
bCPb3XbiuuvwX/rK2dEPsvdNV7o+IlZdNvqGetBPAmvb71B//AcbPvsnpmzBBNvO
QTNxZmO2ehsSEVwc62/vn3DdAx8XS0Bt0tBnSCoWylAm7QLw5voYR6fnM8I+0Ls/
0b1erS4td/amlPfT/FLYFyGyetK9H2YR4c2ADghbhryycsG3/jOd4nPMHsRvggrh
zy9M1iVJ/lDXj6LaNJEW3chPiCafnCr9vWdKtPtWGIBpTCdFHK342sNTfW108B3e
90nTJdOfPH24dazTNpni17IPbpsO2nYtXB/bZjpzZB/yaqJt2ohgoP0G8XNIjI2U
7aYlABIl3sU+Qi0N7E9y6I62ahtT3UzWGvjTBtUeKyFlG7CCAFMpxQyvSCZlKtXA
Uk0NOQxff2AjpadYgpa3421lt1Xrx5XXZW8n9M5m7XTc0DFmP+9jIaiQJPr+6umQ
nCjB2OBHWSAxDInAt8VaChW5KruioQbtNJEz2oT8cTT7qXtzYIhzPaK1reuSI1Qd
UtGWmO30Xeq3OK0HEWu1b+Nvv9jXxUNLJ5vvuv1NvMoDvqvw+dM+kzOPz4fumXYo
FqfbsYheyje/zYSRyrLOphDu9x0bVMgMEWZORysSFjOZHl03IoLW13GX9ouGVRI5
BQNIhCPukzmzD16vLkIqJT24MnOS8wI/P4BQ0k9Cx9pHutPzgJuOUw4V0fbH13S+
NUXOxYdEoorKIl2eFoP9n+lDnOHRVPnBdK8F8aDn468VpQWljxboZF9/GKF54KCt
OLZh8fnC300644BzTjvGZo8y6c8AQLD7jkggatA5FKt18Xfhw5mW0dfiu6tzC3cV
rASnEeiLhmGUwGadR3D8ctaCvhL2G6UVeQnp2UMzkCpDADpzKYhnPrECjCRDScK3
2ZVyJKun+0IJuWsbyLyf3AqaHYm5Xozv7r+/TPTod7hh5Fb+LEpVuGw1YnUDkRc+
miGgqvaFCTLn54WBh/2g3MjiqWk3lfQbvrsrbyZvOERF4yr3BRA8Dt3XpLDM0QJj
PJgfxwfqFGv1c+YD7LjROQdSBy0D3juwOJ9ivoO/8gTQ1RTsXfhshCjXp56FejLY
Tyt7lYoJQKuYCmAkGa/O3NYkjQjqlqXNZgXgOj60aZt9a9nW+1Serdv1uolttqq8
lpImM/gn++guiqEG+uKeXSABXv1mGo2ULEvtFrSQPWHrm/Ycdyqi+BDV/f/DXGqc
VFz2oPe3JDygQqyEQ8niNSCY2sKaCThcHVxaF8Pnz3+SRgA3dfD/gQniHczL7qub
Q1k9WNEpID3t3azStce2ZwhHJ9dE5HrcOFftRr2UMaNgfhmco2H8GjSXimKjIqx9
jYteL2RrAG1qA4B9FMXSNt4tOWWY+ByrSMt0dL9mnXFWd3mvL/AasNd7eiGEQPz/
+NGwikWwbZcVJjcfnHNHBcaIM1e2yrTXuiDTCrF2uGv9zLVhLZ0shPicMq6r2fCq
GCx2mSsKTpynT+wssiD+S2P886ep+2XGsDl9Ap/bw218yAz90BUtUCnp/nxFzCaS
tQEnDK3fQ7IEPhdiLViKI1kiKtRDw9/4z/rvjPATwZQKgE8FgR8FOQ4Av+l9Z7Y9
MY43mlBY9EsQ9BgvhOJ5gNkEeBlzDpDa8zy8zQ3Zz866NcYL/4jE5QRMRvGqiJvL
B0i0V2Vr03ObEGId0uKE/wux3NgASr0uK8PgA3nAl8HOZrJlxJWIgo2LbzZQ5ELr
32RGm1t0jp3bKPs6AKMo3BjozdpF0BL3eOsLo5sA5rUqtVWh00KmepbI44xE2UiW
QDHcS1GfxB0dcLTrDepHY6Dn0LA+X1fb2bHqIKwGd5ZGCGyb+i82AmL0mL4/0eJZ
qgrhtE5oJkRLhtoHLB9yHCSYOUxAn/VpU5mdHb6KU1f57sudsRnJJI9HudtVByAI
guXuayEdFpv37bMwEDWEqJrv8qGZ+K+L3A7ihklpYBxu7O6JHYtaCch70+cXSsPI
mGZtPuNCB9JeLsjjHgLjcPG5UTVXTrbK6C23OQ0r5b/tz/psTFFZJ/9lOW8SdDM/
mxJTzzVcSw8Z5KxblRY1HpI4+gh9mqBMEUnvlYeXF7Fmj3UuIv+nYO43XPw9K30i
dK+Rvak2xPgEo08PfCIiEiOmpsTMXR4+AER0vk6UCqihuhAP9CTzFgeaRu4NuQnG
dCkO4boJJznRr77mxauFoq5B4269S7DHcd3rqgmqO6cSK6mezpTmA8EdtKwbJbOk
J+hXjLtI9sD91f2fC+gQawhMgX8OiNSVtgi4G2y7MxJ8YKaiZ5WDz0fkup71yt6L
yOwknwYxrV3+bh8Kz5iGEM8milsyQYBfRrjA9RFiEMbQlcsfdXveTzrUnSlGDsUp
xImAt/dh43MLAf0DjJzJC+skpJCzIESKRodD/IRfKL+efwO6OezZlfUMnwolgJMv
exV6T5x04LZFaADM49V+W5+va13nbHaeBX2QTHy/2wvsCcGVx0VUEtdTabsmhyRO
WKu4AYESGXdKD6Gi74cGQrC0eDSksU49XuP5LJO+EOf6i+O9EPfG5lOHnuRpa/1v
M+ALpKIq/Puda+SXPouPVMKRrCG5gesL7gHWvA5TBd27ZEQrLLy2pa7mTPzgmkmO
lrO76+0TIx02+b7dZ/JfeEmfHn6mG6lj9XRc+PWmIAyZzaDfQHWF2TqYPaPgEYXp
ao4k+p1YVdL1DP7dwE2DxFxweB6euA7/t2eEmJi8rfO3qbUMrErug0k4p3rAH3S8
KcJtaazywF578HxjTQAXUB8/cB89hpO3NR9GG9WYEouMZp0iHpcjqvEgyASJ0Rl0
azh+0lOcrlHcZiN4+qyxjqENPGAmSJ3ktKxIzbvPkdYp3wjX5zaSnA6XsvDzLIYA
mERxEnQ5XQhrtwUbRI9p+Ozku8fLadPONv9ANYL7UJx0cf7SI9WF1ktmmRZFvbbt
ha/JOHzYLQV6ZB14Wk5KgH6Ihapd38LrOB7Li/+JyuWjHmRD9/3Khu6boYCZ3g8D
0CipzOn32LjBMXRrbpaFq74mpu2plXgVNWYh6FBHkhdn/Vd683L9NksyGk32fF94
RMEPe5paU8q+QPVIvMJQbSY0Taa0EUNkLXIxPll5zGzus5+HuDbvSa2WljfJDGLe
UL1Q+29u46kk+q/GWGxAqurCF90tgXDmi87asYei026XlVbMSJDdGhhto4KgM0xG
4D9lz7zAM4bAk4IPDgXR5dL1uNYOMUXkDsHKPk5Vk4kTMYhiYlg/5Yw1XoYbwDiT
zsyczyvY/pJYv85LFwHXmEme8HF+wICBl9rUZ0JyR3PVOf7ZpcFhcXZSEfG1Sc08
Yr0DFGMhBSXDEuYpKKwuuPYXn0PQiYw0tkWU1DXXDg+06ZvfO3B27HuzvbPCVQUJ
jenj1Hjl+gAm5dgpnAqHe0ztraWj/MvDYt1auZvfIQ6CeAtvzfxdmZSmb0ZUZR1A
uZLsKXfmdfGlNFIP9PvEgPug8q5CwTp0AgwPAq3StPEbIiAStfQmSvP2EAiA/5vm
+PL1IGFpn6mdvNZQRy+zHBm+1McvKJJmsuT3kLT4yr5eDlopjpua5pOb37ulZCWp
8hdOLy0YsUGGw4XmgEamVsdkBtFejEe/u46AlF2+IIMFDHwfdI37OAEXU3yfMHgy
gB4nKas19JsMeUrs3oiV9jChDaX8qB81JGcwyI9EGsNnZ33COn9Vq7Ae1G0ru41u
3cZVWDIuuMCaN693QmzY2a0iwB+MVeZbWJ8yrz6IV2R4ZAGuMJ8E3+fVgWItBaeP
f0kWLtIwTQT6pnHd2rKGQ0q1iGoCDdZSmbYpsLZOjZTNdbHUUuexgNEaCZkBCpYZ
WuvKAc8wvDbdxsbRW+F1VuU7Nu+Whjt+XV92z51pvQCB4tXfh9RIqdLGxkCVFsNc
n+9hIEcEmshigL2gOya5/clGOVd6Ax7zjSGyOz/nexz+onbOcGOV+5xxuyxVn5cQ
Ti/BXIV3VXq2Cwu7higZDVHDGn1Q9FkY8s4sdVCkFJBFxSgvI53nUTXYNGrfeF7i
JZjtPEpCOCrllyDuJ9PCQd0WjAJjhldNO/bqSez7ZdMJZyJNA+vQt4zSBNPrV46e
Qv2YSo38EBky4WQ+Fmj2uN/G4rMF/laGKmCmuSQ/jnefhruBGqXVV95e90NMOT7t
z18rpa6RBc22D6cUjVimREHIpBBt0ol1ZnXl2EmaQ30KulrPhlJHynqqYLvCNNdR
2QS02jhxSsPo/In5tivL9e5QEy7TELdKCF3gNNnCqbwHasakflkU1u1Id3TTEAsP
RJWjWS0uAwpQiGpaj82H4oyaYOevqy6dUIqVCQ1G5h/MAGm9Uvjo+ohrHG4OG9oV
xQSy+uJVGqXTOclyMHA7buSbu92Rr8KAWxO0JFB7SN+mYadUCrSPTfD7PpLhzciB
Eo3fWSp4H93nnc3umSFxMpl/hZOFNImif1XgRo2p3rfWgh/1dl0e7v2eW8KdbRbW
vFvjx9eM6zAOetPPHJtQL4sT47bIKTId3X77Ns9D4xAm6U/gSMzCR8nWj6efWw8b
txUMST5RADRkL2O+C1cYwwYU+YQnr2GC2vUthQhVkBjF1wSkOEVSxAflB8Fqq08v
em49arYKpmuJDvumdJ+MV/1CCc4XljMaQmPWxGlbht76TH2bYJ6n9zAWUS8E5O3o
sUctN0RTTQ1rxRLsyY6H0RVcA9oiZacyImr4fZ7RVeB4JxWFzN0eFqTQVXhRHMRU
NaPUPHafGAjux1+St6rjo/Hay+PVpaGGuNupgX/XbjzsYTTvOcC44BBh8bXLpyg7
jCHVgvGPbx3qKEVArzkx4FKD6j7ebLxewMfVUQRGnj1YO2LVmEUr3u85amTcokqK
AhYRFZffWhlYufVYpRjkBlHRsYIY2sbs4bAoTh7V8jLK2zf50W76Xr7kc1F/qu29
fTlGmwaUCIZ3YGyyCyFEFmHSH8HWfgwL0wP9m0OvJnGfFiDvZHfK6OZcsi/iux+r
iY0D5tYmgc9NeBmudLJpH07Z0qbIvnKDXG5AD+pzT6aVLtaVB+cM3ZL/DcfH88Hz
b7hHxYgsKoe2kMIRrtdAwxyKfFdIT+zyqsskDx8HLDh/f+q1MQPblHC31GPJieCT
OIzZOLuS6D3huWtPzR3ufoXEl9BLpI0yAYtIJ4U5UjBw+tRx75aO+uNQd206nlqc
3AR6PLeTYm1+z7LFC8fodbNkjKDMHPYzcqEU/NMROIZf04ocLkWIWo/DeCeYXrGX
3AQ01PCNLCeJ7Dm4gWmtbyMokZ4GB3n7/dWEIXXam72PgdOvgRuZIASZ8yOObGFF
O1QLuFWZUq0/XJ9SUV8xUklNAdTG2/vpY6u5+IrUXf+phyp3zkOoRcBTIw5s6drk
BwFkAQ1UUYsu64nULHew0BMX7DgWO8e2+dDqJ0Owi3tLxcmSp23+FLDOakQMHOby
3VNz6BPonnnYQw40BpC1Ow==
`pragma protect end_protected
