// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:38 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RS8JZtSvzSv41Vs25Dzm6+oHHJrULHkG+oDz+rDqrLEdOVNsmn/SoN3Jati+iwf3
Mip8CNemceypoTgBB33fvF9YcButBTT2vuGB5m/goyRv06DNAhOLf4v67G9TlDR/
dh0Wi2RCawDGQ9tTOEvYSX4to2ae9QwpOGGM1WXb/lQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15696)
fKz/5ZzxB6iflwDwxPZHDT7FQtXKWLNhA7KESqDGRzlsp/iFSTOP0oTRNHonbJRQ
FvougmJWpcQl8Rm1vekZVwX+tlYqiMXfTvhxTSxzJq+72SrIptJp6ssjynvf/lVX
Rg50zaz/04hcQDp8XGpuGfsBLFMQ1w8XapxA1ggJCp9G/vYko1rCAFx3BxWAyD1C
t/FLWm9X+AzUxbWG1mjyN6hJVOoiIF4egTkaYrwAka6wj1SETRgWPBvWhkDDB8oY
JDcAea1VNcyQ1pxZW1GXdPYSVCcOyHopSOklSVwiql85OQ5TXpYe8gk1xBT/WUUD
t466wPzLHHNN7V2aSQM824HYcUmCUwK1f4lmrGHJYtOtE9rURK70TDr5Puuj1H3z
sbaM1jHIKlXxqLDwu/d5DOIEWVfwkLwDd7rU5g0P3W3N/9NQwcp781P3zHGClmQk
7knvtuFwCraF0kIdUhv+YRzPlJXt3xUv7B0R/RsDaYfEb6/Z7bhZFxMMsDVTpBBw
CZ6AJsbMkXpvhQISM9ym2oeVfqNpJqWuaov3hm6zhslFJLUcfbUZz1l9CWxpWczt
ca2TowPUv6vwLfvjwGkQ5cDewqx1J0gIfW7rX4RL662YFEFqEuya4faFzgrc7olL
rRolt/wA0lGMIw/xdGrLnYZX9WgDCHJZThoNZfxe8tq12rkIhPAduLzQHnyr9lWE
kgDfUgc+tFGi7ELTyrJO1ssHLYuq7GKZm1h69xKOXMxPWyMxJnbBtMUJi5FlyLHK
lKdE9UcUBF5IJ7MbB/AXuKbAqCpb1tnaLdtcMwi31yb+g2KNyoggfhTswCyecGkZ
3wS2jxiHgASKjm5jqoRsTJhfhNEUyiAN2S+DeAIptOZhazefq5Ad/zoTILLkG8WG
vN4NY7+tUoFeAGgqfaaKiPvrR7BkBZgm2YrVyi92Ktz1tsGVrBvfJGI0UCO4WuAo
knZj9cnEUagRGgukeOMtZ222g0TeCWc+Oz8XvBfjZ5k2l+H/jHO6QCbfvdGpMk90
J+M3z2oUqH3isQAiSEYK/zF5s9GHKU+o8kBlYakFN3koafCE5LQPUggUuOtBgQZu
U7rskkzAJ/sO8Ix7EVvxNs7K6iLX9RiaVgAfKaBCuQ0JZaR9FenBnmotZ38UqL6P
RsfASq3ka/NXQ4EsbKv8ynKxwuekQict/4bCNZao/u9seJWmivbSAHrxrKX0jNR2
SpMnzdG/ohKnupudYno0FGe7rldTkbBDenXG4LazpnyChXtFAcLcXG2TbuQeVdad
WWH3hXzwExQyf2fNVgay1FD1sl+CarVorKnvQyxrCZOL+ycOww4z+s3iZ/NvQJHD
Zu9YiPwBwwQiuXdrt6K2gyTdswk6hak9d2/d7Amq4eRpiGtdrpaJ/aUNtfO2jdoI
Ch/W6dy2oPinIzVUXMoUOl8has3IwejPOwup7UkGI+NU0kU/gFEh99uePlFoqhKn
Ppuyvdnyc26F/QnLTPEoEydVT6uUrX6XjpnsN+bTSGPLjTEwzLnkS8vAcHe9EkqD
aenydjOZih3CeP7Ez3+gUUiaHw7ZJMu0lJdbM+MtdIeXpO+ZpOOqBz3LjVuYUlMl
CvPX/wp+/y9I3mfxr7elQBjP3TwUPR1XyHECG3IWQznYCr7wntWVjM3JxCDcnVq/
hGLg1EAA2etS8OCG2AMSxfLSe2CtC5MH1y7zH8TRL5WJZ0MddP+qJb5ViWzb+raM
4PzjKQ2JgmTaNp+tPGKN4c8oSlg4/Z09P292QLC0ymSq9xye6ktR3gLcVWmuqEVy
xvltrASrHGtL25Sa5IIkV26+2HO2Er835GjtBf63TpZqQ7VQdc0Ta/8qr6cbjbeQ
zsvakWhRDEtWogLUgoMiridBoE89zNEZQX6V/JtprkUf9Kpj5/pODcuQA/SJomUA
IjLSK+va/94DmrvdAqcNqwmAPIinF72PXa2ZVigLwgtM1BhSQAgbMbuaL5XUJdU/
vjbx+8WE+MmMjN/uJzCZIpTcKYVFzRxw/1CzsMhYuAUWS9TabIBRCbDK/2fdR+es
aM2sGY55/BuJiHxEJHNTjGVhsInFgZXQTk0zqf3adR2iR9u28lycPx+VNuZ+csIC
xuv7HiFAkzmSzv8DRRic/MeXrKbIQIfUomFRWdHbjoajeUB4MOWuQYUKAdz6AIWA
S1aC2+fIpi7OnlzK7+nbZ6EvUBM3+KfCHrait8wo22GRBfOgb59qB2Sb3S5jDulC
6wDU9lgFKRbwakdxbkXWXv2NY3FA1ZUWZMDVZKbyvvK4dkSDdA5DGEp8S56WkpAz
qo+IILJ7naSOBtXXKvHKwcOTIePWUMWnyzbJ127mMASgtmJJJZAPwRwNs6Jxmyky
75RS9EHg7NGM1lzbn0Ymjq0X0HC/XfYlTwRZBvxx/EA02hNH5WgNpxbRXS3gpLqr
Xyz4ObvlvZGwndr0ZHMxxEoEvOwCbmDbSQR7dY8qGJig4obBH/zXvEFN/XtrIXxP
WmoOyak5jLLsVcY/pdNgMaFtA6bVMypqt00SzABgW9HebUmS4At8qyILJcVV+3y9
fCwK/VUTfki/qL4y/b7+vnYtE9heG34HVpOrBbWmwTRD0NhlhscJZhRNh0h7xCSv
KUiluGFX5LrCxydGbM2Xy1HFYMAHU4vR4KVZGWUxe2EKMv6SuHKGZbl69/hSb3Lj
O/DRRoWgpPSzVThKd+mHbTW9iOIjtpjK+HU8XJgudqmAEZP2JEm4gmLcVggHxBBn
L2WR7O83TUM9zlI4/SRfu/Zk6oKqj+NL5h+iakqR2HOcwI1+odRbKhzLqWQJhUSo
MwAkFG4VQT0JwzZ5EtioF0fpNVwBdJyzHhpl+PQC3gViKDBAjBOmhLdWwCv926N+
QYmzMpr5qrcxzLPfzWZ8+6xjY4Klu3dg/cDV1jrpwdl4viWzbWL9jrJJshssXip4
HHyJmiKeza/4K0cW2H6pRS9WbbLqHdZKXedewonq9VatMkNnppGLHHTu77Opkr3K
bbEiTMzoH5MBIm4BBWniD6OidNSiIfWSBuDre63rqlRSlT4EipVhr1tHdJL0QYa0
nQL8M7B2QsaOAjrIhFNPcqEKEm8tIfWlXGI7+2EsQuno2rtYAklOk28TDNbvFIYR
BRWagd5j82I3bD6sBNaGWNvf7M4meFB0eGLrmq2qTtXsLB+8EjpdWSoItUTW14P1
MvFEW8g6FKIdwTsM+YDkNHovCqkRCuV8nqSYU++qcnFxlLnX24mgm+HyyohPJfyI
ba/BZoobHcNfkn7BiR7XcLXMFveePz/rVyUTSsVLORnQZ33wm96iXolQ62OJpBYj
Uma5Y99XQ9Qyspt3fTtv2C1By91pp2F/2BzCWJQmRl6AWCOxkmWmsIFDpRLgh5v9
aIZsrMyKADkw3vnEvcFjzzPoeE72DNcGCx7u4u9v7gYb4WOAmuWCuRrzMFUdeMcu
FELDFhgOgQusZUg+airYcunjPc/X3hnvssvhsCVYuj0/0R3UpSI0khY1LHjCqz2x
ScbKzsJVcD940tfAPKjG3L40exODWe9rE6/bUmekyYAhNDZS1o0LOE2fPdBrCZeu
jcPPGq2pLgIvDVjW7cEwAYs4EYQlOmmC7OEatgLglNzL8p7WaSyWO+qW54O6Xz4s
6+UOaqOW/KefDJnHGq8UcvZMKWCYJLtKePn85tZ7kuoCUgd0PJmJr0mwYGiRC/3n
/ONtPp5aewkUy4lC5UoNk5S6lm97OC4wenOSm/8n1lyNHQLBic5NnDn087pXpCrI
UF4IfOEfN80MWxo+VLpAeaLHsTKgZQu4/NRE3IQwmkw1pDZC4oQw8RAT7LqJfgdF
usFWfj6gJ865CQSnZK4ir2mAt8RgPJ+WDZ63n8i4hnIN+gq8xWtU3fYUKq4bsdNs
J1/v3sQrqAynorVF7I+qUzntZ9etTAGGtmVJ5CcRXo8QNQ6zHHFDd0L0gyjIth6o
MFTkXwdCMKyNRwoy7pLhJHL8C302f9nqcYcmlRG2pwJzjO6BuRKVVzTDmUi4PUB2
3/t9tYH/0lGr5wgFOT4LQo0L3F2ml70qy+JT1tOZTDg08oY+VcQlwuT6YZpzZ2Ya
ybWZJWnldHIDu/rkec+2YWqxlrcu6j7D8H7ie1AnrjdW9Tnbh0IG70ZAS/LjTZHW
vQ/zOyNv82N9emf3Mev3syO4ovewDt64/GmDiai7s9LZpUBsyQ/K6W2qYyI4BF5t
Ri2Qv5vlryLSE/H9ZtXe0aMvB1BNdMMqiZct0h1XqIoZz7098McI84o1xEyyBQ8C
iYAD9r1a89sqGuMAaqygBRwZkf6nHKg+q51Gqmin9JyXVD8lvEdwVXqSoI8pM+au
1DOzMwNnGJZh5FwfIa4WwlQSovRHtL2BtBKZn0MFRzB7cVGmx0zusb4a++sSoamD
Zf8alCWo1BQv/qjfB+mPOXv3CFbp4T1puy6o6Uq/YdzB07UFraKWw6o9sy3hLVBz
yt/9R6oWI30NDLVPzugSsJMBNJ6LQrDjO24eswIU87Mg9X+VM8s2NHyHcRkjse9z
WY50ebVfDwiLRIqZrm45gNbNELBhKWM+0CrDpw05OWiGWlEB255ld7vWH6hJ7ULW
PzPZfF192pd/08qUVxfr7ELQBR4ucEUT1D298blIzghbbO1OmCYy9Ui0sa+FWp+5
wgeKJXKvw97uX3CGPv9R9AZkYozi/9I+O4Vyjp3MJLC0oSwRjPPjdW2zv5UTk0bM
/yjk8h/dve1q6rbBEHGHaMYCMwg2Fzr67nfLj38z8KlJH7aqwihd1qZMoKmsCVL/
NBL91SxiOzhbe7JfImmDsM38Uu8cFMuyhzYAyzBTExk8Q/vkFAWWqawOZQJ2Jfeb
pdXSqODSFF5OLVrteXsmbwQnFFCi0sH84KxhgWD8QUq1/2Nn97OywzuhLzefHSmR
H1G8f+fBCymq8N/nvajz+wZFFQ04zXDOONDdPh4s1uxkDWp5waoCqVOZnFISe4Wv
Z1D0cSl8Y9x7DdwxXP5TL04mY35rawCegZHda8oqIhIwVv59sIVJPIs7YollaoQC
1elfmvd20bvpV39DR59tzZxwJ5Fa43tZAPnePLGrQUQA/Tqu0fPj4iczJn5CCZgX
TfFlCwm4LuPK0WI0EpGe77dBGB3pc23oDJC38NwUmze+n7oJc3sPWoRV48r0Q95I
kyejQUVMBRA9m8wyaNHC93wEbpyciaUlDsHCCrhdIiYO2EuqR0GtvfM/QRec5hzq
9oiAE2Hp/auJWcA7zv3DBDa2p04GD/VHrVHngv3aNoWzUTN2pRILq0390f5iz7TT
xIMdkEO48jDtP6qgitLYpC+jan/RRfGX3KA38e7RyZABkPaweYhiMbz69hO/5u9V
sV4iSbKj8qDnmqoV5ok/2AZ6d2OEZAo6El2kSbh30uRwoGOBH7MaEqd4FXVaE2Vr
PZSAAQi8zbx9VZ9L4ag6mKjDWU5e8PuXhr/hDhpC7/OBdoSuN23JkQvDQTyoqIgF
xC2Be1Y1dQIlNTW7v27SlqqLgrfgoMMBoC7f9kUznQEsgG4JqthFnC5eW6Sn0gVK
kDq4h2PU8aaQP+GmXvAIjJxs02WuijEGy8PxJ0aK4MiKaTZpm5BJ4C6IKOoUmd5H
YRjEajYwjxRe3Ve/QrUCETm3bRyzYxqBca1ETYfUv7tbpx4kM1fColnoDltKI+JD
8Mn9GfveuGWvflqXfzYer6Obu556pxcTt5MYksSvivwNYfDIGiTSkcRVjf+eqpi3
1w1fW9uJoAsgxoqqT+9og3ov6r748n9fivvBo8hKjk4Z3bt7O5Lo1ILRuMxYvDpS
mcIo5WAk38FJqombbZKSlweydONzkZ10NUqqrxxqtF1p1kP30FE3TnpOo5+mBbzI
G3XeBHEuaf+ichAmGoITeiX7D3wjlu3+D4zWOZ5PllAdFQs1YgFA2Zw0mF+4nJyk
6P99jvTFQFM6vTJS1bKuHRzhBy5f9HTfj6A1Tj7vTzErralo8KZztEapf2dgAzy0
lWN+Ej8IIe52+JDNehBEAfxxtWlyCIzJ4f9iHoIb9BJ6sVaWu2ygGigc69AbHGKk
KbU2PN40gfPf2NuBSDT7xYO9RIZOPSps9DdAzFbu6KMyQH9Pe7sccHJBb4F3LqPg
jMwIvYLv7ZAHKGj6rZlmrN4YX2b3pEfm73xzmqHkwTZxNn8k7lC1wbVS/+TLrtgF
duTzMSCOkGjISTvVR8MCB/bxr6Vi19oP7KE1rRuFBpRe6YskRBGPv/Xk8xoAAk6E
xqsGdZbgXuIYGmRNknokH/GbWkIk3f6dNycs9JXyqweXmxxLI1kNakpDQmhLoCTK
/VeZoRsXci0X0bxo5MlvGqmJJMbnFjcuxfzQwj9XBr0XkcXmcOITuPrGG+EpD8jU
DuXP5XIkYOkhupcFLcdSE28gwyyCxkl1sBpGt9Fykb5z4JhARlPqkjEbhCz03Gxx
75lUDG9T2/UPptk5LQHjBUdkItiRdYEnu/wp0LNey7lWQFjtfKN/RuSW/6VAgKn0
Q56g20RwJcW3/f+8spVv+jtJSO/9V00wStre0zRtSl07qn8M+3KeH3gPBp4BYBYJ
G7LVNMJptZ7YYGMvvan220rgfsm22Q68bcUX4X57JjruX2PNPAfFDmlyZR4EquDH
gitOM5ojZR8WfYMFgbBi9+wdlbZ6vu9fpO3AEf1zN+bHl6+ZmfECLV8dYpqZcDS0
qL+wzIH/IDpxg6ZWa081Qv9bKTmvJFI44cC/b5F3CmJ5yz9zY7GhuOFKMiX3EFTH
oicAAKc8Rda3w4ebUmJ4K4JNCmT6W8swk9zO5YL1UNPMNVNSsq97K9bK+BSLzLBU
FUqs+AyQdfN1ymCzx8hSkTmgKl+/gF+lCHFhZty1aLQcwFDlvnBqZe+pat7/O66w
BKUFvl1tgHhYRhJdSwNL6ennu1RKPFZrwBHVH8W4/GaL51QgN66Z0nX4zykojAQE
2Ln5d1s+OKvvINGa1D7vKvxGhVYzbLLdrf8p2jFpzF70y4o6qqQ/HyfOLx00IYUv
HcZUMdtY3nu69JKS6qYnN9+EBjDIlZfeb6dKIFkPbryMo/qhc4XkfXFcsJyQ78Ef
7uQfHFCEM3mzLN056+xYT0Oeo4ikzhOU5WJlBsPRGbUz6bll06w8gg/0VMJrBEL4
mKRUxJ1lK8H8fv9RfgmQtJxS946zgdgmvbf/q+jmJOooswnr59Cop//cNvoxwH9d
/SuZAuARdd6qPWY8ZtqD/G6n64r6pVx+0d5xsREKjJsUd8WwgOBEi5CvjyTnLPc3
uNrJDL/MSVp7rEdFj2HFWu7V9L9cCyxvOLeIE93Y8GrcYBVBj7exvE2XfrKT5yJ0
eU7z+dvaR6BzOvQOnJKEGhRVUm9xnlxNZjM41DTvLCWKJyBwtlKFPUgcupufSL1p
nn/O8J23c/pZx6cme/GMAQ11LwiB30xrtAbBx+8bEzWZ5efDF2JzGlw5IYfLvkos
hJE561wwzty4SA6jdRpY00xi7DlkUpVzd61k91wWg9oo7mHZ6mx0nZZ0erpLaSmc
hFXLcDl2n8uAu1OZwzyFWjIWEJgI5BVuJvOAgl/eGZCqn22uCgmOWqOj505uaA6J
XLuSC7Nnsc8wW6NnTHFcVqLHRWWwn/adA/oG2qwpeIz282bnUxpY3Eg4ThPcnwGX
43WKjsK5EaAoJo/akryC3pCoSvxfXd2JWY766KtqYYz0V28KKd0JK0NNu8amtCtc
zZFoYDRlh+p5n/qo2DXmkG78ImD2S9ukUrq5Izg3CKgOpt+R+IZdtqCYaf5xfq4P
fW1ZoRhZQRHXQx8RiOVL7uoPcWA1awVA6NF1seApiQUoDFY73qjZuz+CxR1RHsr/
VLByUmW5U/pEstq4MTIkPEqRSU49lbAtLXDmSq97ojbBYu29gisLwYQ+iirO1rDR
4WbQMmNEMXfe5um8qEsULWqlJb69DhE7pry0ce12cEWYVW6PmylGqrA/EVjSmn+i
u9iAI4vokpNDwcLs7aEpcRL8bXmn1VOvYAkDP+2Un+q5mxu2QHThECAWduiAc/pm
xSZ6fbnLAaSBV4c2orqcWqZQpTUxQPeje+uwV2pYf9SuXAHSj91U1unpjjgbi0U8
ZJftFuPsAA85Z6k7fjiPQ4jECjbiD/+0UypXn0kk1zYzNyJge8bPqaABKBXCJxZO
4ovCNzas/4uvQdpJ9e3qBX9VyU/MSHKEBdO5fMKw6bUVCngPCx1es2GrdNCr4qYL
O7zYdDNeic7ldDIVBkimpNdBOCwTq7elAfkKnaPBZ4DPpnXvBPU4uNvKz3GgeYNF
3NKCKNWVsKYoJDntLbx8JqtWrAaFv5tEE5OoXd3ESbWWDFYmXUDgj+fvei7eV4S1
khrBCQDjDrfN1ej7CB4EiE5QbdfqGP74RVeKMA0T/qmo03VnGxLThtIoZNu++Dbf
DIbBm7bkQVd36JHz7FOV+bq8Hd700GhPMYKK5Ehsb8g5yD5a2npoQy5NBFclxt/3
v7UXt5e82du8QzeaFDAvskWxg6qP4bZi/tH3IUjOmtHEXk8Zq+s0CoAgKKO+ripZ
XnvQmrwfJxbBDxxohQBUYRx9CrnxjU6Rn8VnoIFUDiqn3e2Yl7gCznkshwwp2fik
DKqjyPgd7Kv8hqKpbpl9nP5mxc6K9JhR5l4Ilv4JAGG76IXZ3LO2zigUNhRvEy5l
Wjn2rOxCz6XTTx5nf2/AHAHIQWC8vOsUbz34hAemas1W9EG6vDH2mgnNFaKYCgLP
oJRw9Ayk3AKtjCjNXQKdcceuBua6B56OZMS9XIaY3FMm1AwATWJEruBaHUJimwXu
DkAfrynaeyIJZxxbJ1bSF7hBqC55YqwTwsAOO+h/thGgtBti9skhFk10PQq1HkPU
voHPrPgsYNQzHP+SgowQw8ji3cAj8rfgTuiyJ2fsCUv1OO0BT2yTYMpgKKxZtNje
6bDeheYx1hQVK9vi+hUcoN4AhoXJIce9KY/aMZJhwHHXyr1SSyzAkSkMg7yuBoWV
5xvEgTTtjc/EtgdVEZZ7XGrq6nE81wqPRSHJblLyOE6gT0R0/05rEwcTh9ZkGJGV
vR8bjAvGUT1CXMt7+KO/JJgDhP45luIeP9Q0PriiUt0OnKgVDJl8fI8wEk+XlC5x
2TI/WaR9nqHXPlUlMyDaa+FjDwxvdCEylRTKvXf0yD+WJWKcjEnqxBe6DUts7WZZ
5mGKRR7bHF9KfIA3B9Ruqm52bcQNMLNzWjepzwMLBO3ntW6w83BX62+yykcNpp+4
ys7d5o9eJMxNOQuLN0SSTbCvPO/DKtc8KLAt8HE3B0TVRUFTqOs9hxcpzF+uDgS1
VTtawqWgQnW3sbl4zWjbRlzp4VMnLbAkvR9Slzye6cQiGDe7+QjH048e4mGVz56d
5ZRny6peeuxPSPbKukXr/rFKYKxAQtSF/ebh5h0SJAye9tMNmRZU4Qdzt/WicWA3
17oRECWu9prfXQWvag26hR2mAVT+qlZWAYXfivtBx5SXEuA0BC2lkuzcalWDpx3k
Y471UPDnICMKW8cpTQDZ7ObhclCpp/DBKd/Qne/gc8xKC1FQ7KUG78TofRJIClTD
aPDeJ0ihKusqsqMl+elKOZnHn4oCeoYk1O1s0LMcfqFzuB9JuML+n1rSrXEMYo9K
/8fUmqpkEnkCimn5lXapFL5np/rNbt9zyrkkiDA0NiDf6oj+AOaIL4V4reHzt0IK
7vDRohciuAkiX76LitBhux6Be2alFwtuLrAOcNyeEU4WLsOQNCxEoPGI8y4lvMd+
wP8lg5PDxufLHDXeEAhM3njOtm6Oj8cl40XsWuqxhX54BLSrP0+fR8buMoLOS8xR
P3lksufS7hKTlbEYat54DEgLSEdvBcHut5ZQRmqRQDN/Qszyy8QgQAeaeTOTuMkR
A5sL4LU/A/uB2Sa4kj607C/e70JaN931Go82g/VT3+BiSsKY7/P5YCMF61t6oXtF
HH4C0Yg3SKUCaitwzrTNFz7PyghNqbK42ESqLYtswVSa7EOO8KoJxe3b9awL8cm5
15GUNib7uKKZav4DZzHjWPEyYRenKvKrobAsaYzvBuz/vEc6dDqvnoMvaqeTRRYt
k1xCXKwyEdLr4v1/WoBN5+3VqLHo+5zt3sQqxV4B0HYSNes5ASg1ZmVzlcyrqFto
mdPHohkJXUhU9tW3Gin/8Hu+lZNCp2RNZEfEhFP6pKXlqKbU0gEtonJWCkRtBUyn
dSHhx1K7HO9rhhhL6uisIYeZKbe2rQK7hEiIL1yx6So1wFf+Vzbnwruk/y+VUpgg
ol99qEUrXhk9MKRaQHiV8EbbFzKwdk2NpfWT7ImhH7QI078HZPotz632dJkeORzj
q7puniCl6WL1qCM08FaEJXkkhkTAqsHeKzpWWY/Dp882QYdUrkm8TLthHjQfsDhA
8bb/Hj8GTUMGcFwG0CRplt8/P0Lqo6aRk/g9gV/Se0iFoHgJRs+EwChBKywuGaVX
aYZrdGTCDFBd0yuu1KKX2vlcsGk103DZIIZQIPdP1zTA/BZvko1jrqV2sl/9YlfT
JV/DJqaELn5k2GewKeR6NyTaY+eZQ77uXwtaatIp1iHzd3a4gd3nPSh6w5+YMGHo
2n9sgZ2InKXEfxfc7ceZ5DAm5iJQE1YAC/vFoC+9F/KS8VCLoMze4B+EmdKvSGmx
3x/puVpvSuPS6NUVUBEPXmYLK111Kiwg9kAo5f1oWOmv9fexe5iLiKi45w0WVAhv
gliggCVyCIDETNy71q3La5LSINhBWfJNINxrpbuO05V5MZCy2F3RCQf82JM8C36N
r1mUUERXMmPOoIvUCpXEOZzOniE4nEshyWNDIpFO+/Mj9+8IyerFWxdqEHLEw2an
Y/h6ozRUMkO1ax5gQJet984RV+ZeOiXG5mtzCIXJIcQX6KNnvhh2vS66Qw7Px9al
zeTwFkIrsqkgZUM+A15pUVpdIHSaUJzW0ODr1TjbPxSp6b3kwnrA83mYD/9mymvv
EMW6UQBSDyk+R1oSwDwIud8WrDyawRBnkIUhVb5RE1CytheoXsqe+kU86D5JM2un
Za0YotjRpiafXKTlWz6gFNPgVXwuk3qtCvas0nX0XhCQiZ4L/kUelApF8QCPgMKQ
BiQDuFp723XeEDwHFJI69zF7dHur4zav6KcOtkkvGIPKmu5bMyMqq0fndb4SS1wv
wF/MxwzffLMlLr4hCwMIAOzl0K6NbK6ew0HQnmMvsC+SRlHBX8e6NUh3r10PYbLB
eBQ812lbASqhPjNQszzdbCIWqfDpLqW/dNJFGZp8h3pB0IaQ8kYftLx3RlARYn9F
4ywmfWcMnCLkWRrUuwq0bCSUHCsDlZR020bsuoc9Q8tKyzLveowtgIf8cwPdKa2H
WdAenqBZjxYJp1cVYMU6IvvDkb0dSP91SwhZy4SRgFUMnWA8bF7Lm8F889fY3cNc
0LMFgJ5I7DvH+Ry8E+XpZncoelLZMavCXI9pvyWDImbnkZU1/Q40ojxGE/vhP3wh
0VJKpT180eQyqnaKwV2ZEY41eMWrwvYEs18DMCehOfPOS7H8WBRe41gpY+RUhwBr
je9dYNGXgenZsrtfbVf78R7a6srhnNYZlVGJCV6G2sZxUQiNZUjoXRfhvKaEqjbl
jcpLnPuHhhZ/Axactq7nGG/qlrR70nbmuFTZUJa88S9SI7jJsF21SXeZXOuWDGEd
IqE0/z46G4N6SAZrmGuwhW5v/zj1m5LH1qSrPe1P5H0pc3vGYdAFT1dxbAFw05t3
Mecsw+gAXjWzx8uohpxIC1XKrOfFBT5zXGZi3+BFnN3B9CSZrXaKUnWchgxrCxhc
OesbeYLgtQj4u77/Y0d2PuUTwIBdXIcyVXTI8YM44lQhRuXky4lCY7YIXhFHrpG4
XUzDb3wH/6DdeL5royzCIS6plF32T9D8uQ0+OJ+EejKwmiE7TRponxr3z3NsliEv
eBx7GwBB9T1tk5666MiiDLi0Fk8MsKrttk1rKMY3IgIqHz4uLgrtCaHSGZnYPVVz
RezRxGPGmGwzQkU2slqGibXtTTqnc/txaeNHm5b6y7tZ/HA1pXrwn/I+xj8nF3/v
d/NWLCKdVokDnFBy7M2hMEqiV155wGvGZ4tLHQADda0xOMWtv11CQlkNQSW81rhX
lge+FSQawRzmj6Hw1pzFjKT9lcTadFDb+m8BG8J+WQfMV5Em5Z1P+ELg4YlXMcyD
KUGQXOCpALYr8uN9szPuVVJaNettHMB63mb7Ih4gMFjdMhUaiI16Tf8fmcsv9og8
NE0e035sRK6zFGgM/sp2JbhIJy651t4ZSpn6ssUg3wjMyILNNn2cg4qNMvJ2FBsJ
QM0Xn+PyLJyo4SlIPp2A+hyRlqCVR5EdWPhObmnc4FbLIuHbr4utEptVO0Q3zSUo
dkoaXgEIbUDt+Zkbc/rKeDu6R01G0pWgfROXBSZ7E4amoq6RwjrsTFpyJe935tna
sSmJ5El7HVIMxfW7+yFOICiRQBrUo80NkfTfvyFK3sMpAnISNsxnPg75D0vdlUMA
JUijlcnMubwyFTSQacoR0m1WWzU/cfgwpr4ArBvUZE3So3KBIIzCdQy6FoebOA2C
Asi43klToK8kdIKKTHUColGjCkoelLp4aonAMIvgGStF0BB/mHxC+o6lB85BxRvz
4QnOLp5dF9Zdkjw43brokg6k47y9WnK/BM6ysDpRPezbzLr/AnnVYDHuTrEskezu
XiQPBc5k70fzhisJKAaUD8sJlS+sJ/LRPTDRXpimh67JV9K2DaX2oxCwwMpvrX6K
sMmQyEkAoQmjBaYIicMNIJz3RxckLrjb8X0dPvLEHl2Q6/2O5/edIL3YQyH02l8i
PadLRtzrVHWazpPQyHLB7JqHLigw3CscG1+L2caVGRYG6sxcLMkT4ywgBEPo4IMW
jjuaMvj2cQzRZCRPZR3g56zr0ZzFxuzWoXCSXsw6jZX11ncLijhhiSoA5VnD+wcF
IFgfxK1eGYLuHpauvXysdUuCoVGMv0hArCOzRFVE3BfSS/prAS6UPUsv5F4KCi7l
iZnk3l0N9vmBA5p5Ekfe1pJYzKIZhASV3Wa3VF+1jE+vB+zBx7ESoWWvx4LvSkFW
yX1tslCcMOSLxaMIrYtzQ2qbvmn+BT2vnu6y5c7z3Rdk+mkGNPFc298EUQ2AJJMA
3tmKgtHpOsGXTC59rk8XctC1d3A8u6ecTjZ1rq6x79ODZVF8wQsDctgDVayXVXnR
Bi62tSI/2FGNf2gYqf+QacXvTjt4rfgPxZWZHdEdCAIuiRI3cM8aQK2AGVtyXfHe
QdZDj4zvyS7gwKfEkWF7c8RHlKx8FJZA+zogVzIthJQIU3f5pE8nmnQr5iVm35Gt
WVXlLhRegq+394gPwg3NndNZvhZX0NVn6IPh6Lxf2iL5VMW1QZUbOxzzA9ETsjcK
WxFrxiswJIMgv4PRpaIRVJaD9YuaAIDwFco+lix8myzZONgfUyJ8Dx93vjCeO5IC
UO7RturMMIrZRaKbb3gSPDdKYouO+5RI04fCLKBl+K4wS6+QazPO3uHHevOrwaph
gPIijOU/TnrQhjyXWsz0zPV5KoCq8FBrFT/U3UKRClVJjPdBslfR0WetthCUv3v9
hd1C/niJuTh49j7+VLXBYnZ+OQZ/AHcIIwbJISqOHhPNpvaXyrlvPUz8QArwFYql
9KceIejgtj2FzMwwtkML82dh0urfIrQ0lmuxDaCxpIltwDxYQFDvXMAQg76/qz9u
TeeCtr+zPYRX0ZpgtLQDDxDmWIxLmFnuyLuBXZb/o3fM6dN0LY9ZZ7yDHgnZwjcj
vUlBrxARSkgBAqrCjqaxmRMt3aij9Up2ScWeoX1lydfAPbopzIY84183z6N6Cx90
mo1FHtVNn5BYlrq7H/4ETsFm8pm2UVgT2TtdnOrG2xTXP4Y2wY6fRKlNn+ckM9yZ
xm3OmDlkKyRss+2rjtlBf0+WyavKK7L6GHNOD7AihPy5Wh26aGWzgcstti3EJslQ
Z3ESeG05wgLRNZfFUokRned5h1PL6/QlXfFMGzZe47ywapGKnDFoYQYTnLLYENIB
mq+BVem/YRfhG1jr+DXOswC5Mj0BRM23f6PlrptDzjtNrfO0QNs1pvqGJD6EWb6r
fS5bVLMvzzDYnqWlOxvRetE3E2rA9ane6VhkzVFw2wU5h1f1OTIqgY7D6EdIW+Fh
UXCw7+WQa+GSdcLVR73n1CRgcYJquPcxjmgrqwuoqIKaQzagVReTr3b+dR+StRp2
PszhOPf6fd+MxGkQ2cdX1bA7rCp4VdYAYVPxY4x1JmkmwmCjhvkjf0n8GrqztpTd
HZB63RLE73A+TUmhYrSQdB0yXeBkgb7c/7NYDrMw33R+TA1IrUaee213C4URf3us
3eUFO157nb87kM6l4iqGBiR9ELt8Md320cwLAv/rjo1RQPJ1qFcin25KZs8FsL8i
SyqlQGzisT1BeTO9GhrhcudGKV4RYwtErWRUIj4IcHJFC0Sl44ibAs7e8qGoojKl
AFd49zAT8Jk2CPqCn7y8ggowXt0t7Cw8Yy5E5wcBNHjY+jb1Oc2Gso0A2tL4B3PO
TdESm7aFDgudrZw2xZmrD4yDiml6gTjlRx4AiCdekdf0xYCUChP9O5HjLSZN1YZA
5KvCGuvjFnj6FXhmyd+KPpF8HgqLrPJdan4BgVDPqIV7VRtgPrG5S9bu2Yd34Kwg
rR9CzbGcGWG/oVGuuZpSKneqGFcUHLeI2GsdejRXLwhWc/sgESWzAZkdCAtVHM0I
pgqNUmaT2dTioCX0XGSX1VEeMxpcv/eBxDa1mUObtyieev7s47G+YrjKsnyqrBBo
uOpt+oua0mhPgmTLbnZWCGRYEoyk0xnz5g26SXM8GciDFVNF73zg2+DNt3hE8lk9
2FqtmMlSIml+2t3ISE6Brmblay+kOFbOh/1iEBVgkpWebk+dk8Gpoyg/WZnu2tiU
hEyh+OzNiAluhxTn1OrcuPNrAb6IVRuL+yQ7BuSxxI+tCvxwhjWeOJcxv0QMSOvY
qgY7EfXosft46Bc9UCXrjs1J4+RkiPyU6yt8I6tdzrIYQA2fWG7XQboerfr22VPX
mBbQ/O7IaRpwSPOpkRjNDYD0SNqg1mICO5ic11k7IzEe4Bm/KNwoT3ul7hp/G4zI
aj3Dr4I7FSziiwftVHOKq3X/uN/DW/Plt8Ola3AOUyWvkVg5yquCMkC86oT8nhyL
1uFE6wOz1iaAj9VWZ9VFOQ/VWyCxF+ixV0C5hZ9hx9/5EUs1roqlyUIVwzfgJ4xD
H+2nij8wHPCH5ocVr/gTqmW6QGci0iIzXvu4y+iPrFgCtmqfmHc9acD9W+1Gs3H1
jZIr/6T5JGDNv8rbcEp754TDGiTINa9uqzLxYYoKjYfuNZIuW2/C1mBHZhuIRP4v
SnFZQef3MqTROmjtROTzqIRmsXojdlXsRzvJELZub3BxzsC/3DTN0AS2ITq2TOQD
Y5fkdUqz01UvqWIeqJInHg7+2bNHsleLTwPugu99feH3biFT8cftIPwvF0U7maZG
GrlKAJOk4K9T+J6SoAfWAF2MmmXLgOSWDoWWMnMrI9UmOTPeyqBCt/HjWC2FlUPO
jUUKnAmzKehfgLfKtZkPex4xMeypmKJU6M05SIexkb4DoPQ9RApa2AudpvWVBDlL
r9T7e9EhvThrgnMHeiBJo//VJS3PPMLgrUa63IyA7USTTOyaYO2pmxvJq911WCUN
s/HoZGjv2NK9hSE6BUDoJ5j5hAL+vUIZhcb0i9X8phWcz6qRudRAel56HmDxD4Eq
F5r1rVsGRmpLFhGRR4WX5jd02indpDCsZrquyTGSaWtWVzO89OmbZIKkJ933nVDt
O4AIZA3VJ0iMNiFDcIUamUZ9wsAwUKjJx6ZDKP0gUxTf6BJBK4/A9udnpTX90Hl2
8KKCY+UOkT2DlBVGI6CN26z7UHozFm0P90uNxsuRZDlBBrzaKyoXEVLdAHeypBcu
r7W8/1bYckiTiTwdEB7fvY8VgOPaHTKWwoy5FgFLrw62CjV0CiXQTIGQJvFw7lAy
ayrRVmtOZ0FkufgGKhoKFn/IjD4EsDOXWzOvwJBpkKV+c8sNhVNhAt6QfjykAXNm
Az36phzja8sGgc+Y2wrOAGdvoTDu0AtBoMUYr34bVq4TaUbWWrpMKeaxbSqlO/Ae
rlTosXGm1NZJYYAq4UOPBt3PEHDpiThI5oFfn4pqyis40gEFsnYc4O2xZBwi9NKL
cxqNl/91+M5fy0FfvtqzWBDeuOzkTiHpmVptJP7iwyntyxI9YoBByBdD3dFV+g6W
ISz6BpVATk/H2flGTunyVLVFRQa7L6SCufbVL7XRJ9EgdkuOufBzp0qPWx5VLIPB
eLXM9Lur5c9YJf4DHRM6Fb7sw7Y3x70NjZ7OUH945NipkEprlC+LKLGozPo/fDL+
ajFtZHsyOzXVKiCGUrNil8TSxaxGR/v9ays5JO+I0W2ijJN1Py/NNNxymrX5Vx6B
afD9QslZdFJaBc1JkBhqASYlpncrz5wHbQJycSzbrlgJfEk/XFGL/ehvNMtRZ2s7
g+CI33bi4fQiTilLKMpMggvjbn9HCzq2vjWlB2EZRtBt1jPbQ41zImOAGmos6mXp
vTERPy+J/l+FL7tZMvGVtSNC+ekw3iXlLRku+teSNvq+F2ELdk3qJfHB7fJw74Mf
NfXrGRYvfOuK/4yGHgWhxiPXkY+5YpR4s7Ckh/RizwKs5zYYKQ6eSWO5c9rWT36r
p//2Yum2Xx214r5sqs4X179qkfgzbJ3iWs2H8rjiQpMIlW7HZ3JUz7vG58JhzsNp
aRv12gF9lpgkFxFcPRQRLkRnj3qeoRBVd4xjJ/Wu1o3h31QIhNIk+bFMmVWIjv3O
HM3bMUSDpQUHF/IW81e+ZyjWh+faPNkVDesSWo7zL7/cWf1rxx96LXsn556rs3Mv
rP9Zn1WoewGtWrkBL/I6p+PSBZBGRdNfPaWo8VKWKBx2AH/qZXi37ZSi+OuRUP6o
gCC4x5k5aYAevBSr34FFhbqR4fRsz7QO9aPD6wzrAcPXeN+I9On9g8pNWVP+mg5C
Lr2vghL82wzI1/A02WjvJ+bigDDLshQ357BiAmQOoC6cT6TpD0E5UuPZXeXSHojn
d2w8rXpmoU0GIYzOmEiiM0Z2MXK4XrHEhmHXCyqn+F6evnrauuE+ES/yRQKwDIf6
Km8n7TzSVLePNA3WdsQN+wylGt5mwBI3gwNsF40c162UG/MTQmNVRZUgkQtWmo/b
3BKgor7J6Qh0ZU9wUfCwBzF620EmvZuKC1Vd2wWLcBPneWCDD1C46cz5RzZpbtum
Ht9erEUkzF5sGO9oXlgsjCpzCeGQwBKueQUO+7vo561bjD+V2j32r2ISkncH5a50
UwXV3eYPgAuMzAFeomeF2i+Fn07UA3HuIkwxfdBykpcPyd94wahW6HknSUTAAhK6
HWs7/Ps2VJHlIr7aY53WypF+1sf2Vg2PuIZqiBDNyPtrjx8W/i+hF2v181zKOzq5
4JD29vbpuhL2JxQ/gZF/OWCjSA8G1IRsU/O+O4ZrDXvf9vnT7Q+V6ccYV6DKr5pb
W6K9lS01kAQzgT+beBesrCRD/9sFGaBtTHz7susALFQUlK4EG0I97Xu0nlfo6MQk
bRHe9bVYotukF2HIfhmPxxaC8pYX2/X7oV9zCng2PLz5mkB7bYadD6OrGY8gHmhZ
b+mAWIcV17I2LryqSyfnntwbQWWKOqvJjrnLIqcJTy7J847MOsceiBOqtuukvr86
EkK0WgjFXEAse2TM2uU5TXQv1KVArc8tm7zvSUi6IPlzEaa+xx3JxpRU4w1zeamv
uaot0d1WulUnS7H4dZNsrmEgvJsvxa8nWmqLctKtu0NRucdK1FBiWhHovMHE5DP4
9gjl5DX2v3BVLvpZQnj3lykjE6DcccJt9uHzgK0Sm8m6MKuaa6D/ip3JnCugU2AB
TNtz3f0KfXpdofxo5YPZStJwO1yzuMWGApadtEnWS4HeVXzghEf/ztvTovszS4g/
HcAkUCK87V8OVzQJXmFB6aNpW3pgzD5hgYvEmL6SlrnPnxLn2AQ+JIppXCt/MJan
1Kbro3DZz7OT+UvqgNhtq0K3oZ4a0nXN7NkA0cjik7s0JIuuLqo6njuoD2vS0Osc
+AXxt4yd4NKZbPkKCgCvnkRaPwJ+ybrj/+SHEqob2RH8lcKEzm5bQNz3wWJVgvmy
H/O8r+RqumdeQEZBVPrilfSmsQT7BgqFo+6xRkqsC0v98gUSm/DkT0SJrAm+5aqY
r2i6i68rFp/yqIKiv9mFKetM46yC7lU/sF6Hlu/zbmSheGOsR5PIXc2Ly7riHXSP
Jj4qmenHwUve2p2cA0lo66swyWPI4lBUXiqkePuESd5yhqPWMTL87x6AaRLJ6HPC
QKms+RgPrgeVjbF6Dfye7A+HEsJ2ZTk+Ni1dW+yeBeK1a1U2unQhLLq+stSmfGls
uGL/xe1ZBsi7cj85qCVZfgHRBPnW8cNp6biwcQ65FnInqGMncmkYfel76rz1H/u4
3vnlodyHze9bLjsC6DGh+f3mHGDkfDYAy4FpA8LCMls1yEy+nWTWM91IEIccodiJ
59fM0rfJ4IiJ1WCLbtxjc0jY11j57iLUn8WNyaJ+qoTdXyeXh32bWsfBScsfOlGz
iatJ9NGiVjOxEiF6FVazs81XPWS+BmXGXlkxzusIw+UV0bQVfhYd1LC4QP3ArJTY
ibsJT4FNL86yIitMY5DyiJYjSeqRJXU8JEa0n+AbN5/S0MeL6S1UM11yDGH/sS1I
hboqmFT0MaRszx2Th2FqLXhGcEriIxCWLkckHQne3rpiPcNEghbVgQbLAuNK2+I8
9Coi2V9lBP4+y9/56suP4ooqBxCtvu6X3S7Qg647wUbiLBA6LdkwXXcoKTVqRsCd
TZIZ3JbKFi/8eIuZKosGMhV5DIV1VAVCT+nMToUVYmWkbVxPC3lfoXziM9P84DZW
IbevZIh3U5ZhH8jU2SZGfnoYYDZbLyMlkx4z5Kz22HwQRnfVl6gTmxnnf8Vg/feR
rG7WUQS3UheMmJa3Pd0dlPAUfW6em19THysKKkohVZzY9GzKroenyspaB8JHhbaG
bDRMkAhfHgao4kNtnjsdlRiSkTL67Q9MZ7gZOLupQjrKOX5Z7bXKppapjZ08gGg1
5ACN+q6fU1Xs7K+axjt9fdIOchehFZAr27o1lYaALiXI6XS/VxZM2/uF1iFog2RP
Uj0glQJSGgsL3f69YOhoR0+iWVHpo3PjwW2v0wgFOHOHdUtxfSuXsJ16CvGFZRJb
mle4E4hiDF2mWKhNNXycJucPAnjBKXIyT3JfTFrvufa2+EF6xcSl6NZ3Z6mPkZLl
kBixoqW8J7rWmz/g7p7GKLUQNau1/GyCF8LGR6CBwZRFxDTRnEIMAmzI4yi+FZLk
lwEbrM6ObOU9TiPKWXUC8dfCU4I/94Ut45Yaf2PCh53BmwSIpXvYsokW2UGgO9sd
l3jRdutI1PWuNYsD5heRdzpbaXt6na4MgkiWVcuq92z05bUZQ9L9vGqB4mvK3wDe
g527i/3YEJazWZ72wkwGxNmxxiBD6+7ivXbBCeh2INlYE7HADw1E72x7GMYZS93/
cRXfUXeHRg706XtyNE05fPM4iRnF8PSFdNrIHB6nv7bH7DYOnl+cP1PuuiGWteaD
gmQipZrbp7nJdnWBObAbi9qeiMw+Bqvd138TNsQmiaL8H2tT6iWLiceCdF+Ji0Ul
sF8Zbf3w8CxCa8MYp46U1hfPfwaPnS3GX26LsNN6a+1wona3UvBHalPU0bqN/yyd
JZoqu/mE75rO3jsqEMRxIvBPWCGzgbIfPx8hCfQOhiKwNupNC58yoB6IrjagYAzJ
N/zkgeIwPiINYyYd9zcx4c6fi1iW6Sf7Uiig6HY2Oc2YExICAHpvTh+tjVP7f2GW
lFWBzwCrEeId0gtjNWvSrS9n1SWqv9Ue8QyCyfovIwhFx3D0KAENX4O3/GLYiJU6
BDry5TGk9L/b6Db7px8dSKob1CmAcPrBpW6X0cN+rwTb7z5ofXwZBdnT4yhKANWk
O3xJ/cXhGKHQdGu7Tr2ORP7u/jScYoxWSA15p7zd/3YneGTLg9MA5TcfPqd/WJBT
mWmelF4ZsrojmlrHg2vM5jnazFz2KaUOqspDfuK0MHG9SoeBoDyH6e6JmIjdzx4c
oqojGuE7h7O+4svE0KA5Eur3GKd13/r7ppMINA+ZUBZfuHsA0IwX4Lhoc6mCCEVa
OV0pZkkobRt1LyM0UiC8A+Lt2aXdAhkWxgkv4sX2LQaahmPNxJZhSL7b8sN98cfp
Zg4rDNOeFkqZUHhTe+9PNlXhQAJcdXimf9eQri9dIXlQXHGTqGxfkR9PwVTzhC5X
8D/zn8u4vEma9TlOU7cScSPd/73k9lXmSCzV8qE+eAi1I7xG2ooRnA9AnM0hAV5b
ogHciy7fjTpPmif/tLJGiZajkBGjCFkeTL00+RPjeAcM+z1KBTx7xok4p7JGJzZ2
GyJot+oTf8PO45jExfj+Oz21G1qhx8OTJuYb1xxSXSPuQZXzCQ5EXhnbC+KyTjGM
w/dYG0DvliCWGUMFmYnDzNyMUGVk2kYltXnfIkjT3bWjgP8SEnKN39zzg6D5QT98
NSipw8M7AC4snDp6oEmSsG/ur4CXqru+bx5LAu244PRHk3fF6agn7jwNEvIKEybu
p0Xf1Pqhcx0wmDXV3ANbIq6OILgm189TxrHDEEkaZ68nPHV61O5fLX4xYVPaq4Cl
CfpN6Gw+mhnbLn3bL0eGlAMJdOVPj+XC/y5rTcfek2KGYn7AG+i5nuxJfYqkVvqS
QDpgsK4Ss5BVEiMLvNNqTU7VWK0IfRSxY6cMeOdjCFR8cFvm+ypk2K9NPel0Rwe6
`pragma protect end_protected
