// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:00 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MyVdebfah6Kn4qJDZCdmvsIIWAuFBo50HjIwn565je9HDBqGzU9BScb66S13qOob
tGGXIsrUP7J+z4sYqg6+GSTN7wAy3FrPJrqSFwRzvoVE/MqJdSM5rnWDx36J6Tw4
tPzbes2n//8c0I6Cl7WCN3LK1GNvCYUrQ5B48PHbEpk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22624)
jcP4H3BwmxaBEdUDYUtKiffw4G1sf5iaRuAe0EoxzNGW1aZ7Vr6DnQWbgDqidpSc
9TrIJg64i+YzhHcsdS3xDwRZtljwrid/q/u0neinHkwJHamb1KDGvtfofK6psbv5
memuBb9r5s4PVdjPMWQY99yQyb0Z37uKcW8akkYUI8Fzi3Qo2WtjD3LWdiQIjqEk
kU84bdiYeyhqy6NMWmsFC9lpfzS+8bqW8RxXVOJMXuAA5ueiBFekU8yK4eoZUR7W
q4xzCKWyDMZr5t0qddM7CxSgNpTNaFIQeYAh7b5zU7l1bPHdJB86LnbHVTdpAX18
nhQop+MDqR8VJzWHfxSeitBRwNqDXiLSEB0lVdUrIwPtpAGZy357onrLdjyNbbrp
U/3W775WoehBsAV0Dg6aR9ZMCQim2Whl0OXqE9mb8SGIIF89fvXVTAhvewnBGALj
zqH1T6WEgyoSsjGd6P9lwieV6WKKws8vnPK2KlFBhkbP4A7l1CvEiZakNQez+7jz
berXTcBLeAvLFUnJVEyfKOYLaLA1AJr2XiumVwCCjHIE4uY4HCYeERDE6K5a3Ilx
XK2VAcLindac8uDZnX9faJk4fEhk9BCtWcAcgluK3UWuuOf5es/iMOkXXbkbyEnT
nZ/NHkb9aaSYqQtBmEv13PvU15Lk7uFQa05ioUqwRsSJQ1B5D8ML+hjb1cwO2Rdw
5ysHWDsSAHf87LLKDj+XZCwNCNrvqf2AZIopBd8FT7ddS9qj1zyltpa9rh+xlMTS
Sq9+mdianSfDR8yehtd4cLRnGESNLsEYEmthgwxjwu2j7r4I6K93tQbrPJ5FKvZ5
TpQ35pdDFmNeSyckvaW7A8lHZloOcuVYaumXmhuqamneZ1wr51sevzixfBn8Nm6S
aAISnCTBqBisfyhMG3TAVtthqpCAfmwB7P+82sSWWqJvHp5Cpco2cw6+HqF4anxO
9iZCIz6PprJ3+gLQnXMA2nIgcADf1/k5xiSJ0hwwGgJAhcwzIYINvZEaPp5T5r1/
jB5RwtpW2EVggXtq0ah9AjA+d10NgbJCKlPWCNDMkXWFIRw9nxlau8vCiOyZujh6
xfL3yeothbE4BolgjvaVD5eImHJ4YZWZdJqubxZthMW5OyzvouP2LEMi9cLFfbXm
W+L3Um7BRZs+FotsFqU7QKQdmH37AlUjuH9HegSIXfu851G7I7Y0kxVj8T2avh5g
qxjqiSiYrLc/AEzIKuu5txh5Z+k1lV4VMzpAvfODQuzFb+i+HsLmaPEz69rSwbH9
TfMQ4GxVob+h8kdrXF6F0NAFwCt//MAiR2tdHZ9nxp9IbclKlWm8BCbuNtCVCmx6
qGMn033xgRvt5JUGc++Ono3qRN6G4VZvavWsxFR4Lm2mGglwA8sm9k8VduSeN0pY
732KHXSVIrk3QmcBglhmKWm1txXIlfntKat+9GC6P1QTQOwZwXb4s7u4jeCTv2E4
JmqQhDq4YPX/6qx+QYfyBYGSyP1Mz3ckQ/OKYWVaWAptJ8WRsSyErjePbiZV6pI/
/TrSQYbq4xsKJBopBJW6bw7w5gMm0GURANBFW1dvsGn5MImaINGkNdrhv+TDMhda
A0HXv/AflCBIBsbsSXA+77hRKBHWPiPoGa++UrttGmLw5LV7tGG0t1CbotYQzu2F
4pgL4oN8Zk6yYyjorU5g0czcGZKg/XRtr3ybbb7+QuyzaaSr4e4qSAwDux8iHHUo
zDrnEIMbLYe37L7pX0t8e2P9N//cqSAEPVIGrrOq4TwlCvLUxAoMWxR9kV9H1vVD
E2agwrfXQ20R9SpPq9V5SK8hVhAyl+WsjdRo+HllD9biu9zrtnlZWAj8s6WbKdTK
81E0uxGbW6b6xIPZZb5SW+KDaSxIyBwxbQgHLKR46JP8sLXTgUGs4dR/NOBKiIJy
uUazw6VeVGz5udjybUAjYSq7RmRdOKSIFC+m0X3BF4xXEmegPqfsW+TMWUhLA19L
VK0D/EZEdj1RIJQHr04ugEDSq16Bxel8nwpLuqdiCTOMJfZv9yAh9JJ8SMeiPLil
1A19kc2D0yN6P+dvzKfeMmOjl6QESDzdlbrwxURM8/JYRAMPzSIv0tiRw0D7R5Dr
g24rLZc4W7O5fkFvpeP+y/9PpxYCY5TgatbdSzutBdPq2YhPwQm9bNbmuPnia2xQ
k6QKqGxl7QOIpOWNI4aJhFCWIr1KgsdcJgNjqzrLh1Pf9zvVJETzplWZuuNuzuLa
Sey2x03pO6+b2DMeYWTaMGhAUD19zPKoVBDFJCcyqUeoR7xuemIq5D7Jr1EfVe4/
NMgewo0Nysw9j6Ci816MTjBkIa5nm99aavmrmkljwfkYrHOwoAJcHnmnAhNWyYp7
mqFYTbVH+yK0SXeB585YQjz1ZEz3VTImmOfBKvpgoEWMPnWwHN8kNMATI0XvYzo4
DJraT+7xZ5HEDOadLBcILvKmUT6wVal8jrEchxlrSc82KN+Ax4QnJdrmvhjRD9GC
ViS4mNekXjCV2IYgUlct6vd+JAubKuwJkCaLKSuwS52fKJ0/cWnYGNOWLsRsyKwf
FL0qb0lRMjMHtemjDxjX2yzjmyJyiHz4eOl7CGDkMKXwh4XElx6/z1H8JEJBnnhP
0AHvFjx5E3A/pJ61e4pNL74d+RWWNAEKMevZ6iIp96TbR136UxInajtHflDpFrFB
VClxWMP6qcP3lu+e9etpqp0gxMnL+c+H4SLkvHf60MYqIwHj7QIXPdLnsDQwHcpe
F1i/XHu/KZ6/yrakoUa3tGKQIxrVQtQ/waLVyTD5IX4msHxYusvXkuaKpuWdZj8A
o9/O5YI2VcpHBu2Mfm7y4IjgM3dgiLPsjM9UaLKTHlPOkR9siSjYjsdWF8IOgYVH
clWMf+XdtKgBhdo8zM2jAgaSExiUS4/0GMG4TuOIgX0YvDMsiiSfHqHJPPs/Ik37
kfP+XdYWNKVe2HeKbyI8F/8nJh3Y+30YCT2wr0F3L3NUzC2o0R/UlIvm05ZxGigv
kAKXTmG80kheS0hTA4zB28fIh7sN1Ef8GYqoU8Do2w0EK/ZDlX7gK+TY4SJKdUkk
3uGL/qg2XIy9TP2yiVt/Rp9VrJyibSIja8mMhGmr9vewMAmQTAoLvRXFfX63CcTe
RUAeSosy6OPz4zLbBLnNG0OeqP481FfKWkj4cHpqB8YgV20by5dItLeZqhHyHVr+
FyhUQ1kvNhqPeFazUjj4NI01SXgDtSQmMy57oxp2x7zIt7hWTtsRGYgRd7T/RlYR
Z+M+HLZuVQsp88ortNGonLXy4hvaNSX6IuqOM7hj4A58D+iq5hbaMsTDLGRXxuOJ
sluE6ax0bpQcdfr+xC4cUuzlKJI+3MzLi8ggKr4EQi2EE3/MMWtGZNJ1ZkidCTqW
IktT0M9HMGWOOe6hHs0pdEQb72fZXA42HlDNegcZOZaEj+6kTewzk2uRzCn2KrI/
NtKMujY3MmltnDTdV6p6WzlS3mHvkpfFjYnlnY/Z+Gf2wkHQvlsH9olWQRXmMPUV
Ku7uCaMjyWJ9SEAWlX6e501xqb6si1Ri4eoFZxkCQo7xEqfpnwaZDkatfZa/iJ4N
IMqA0v0LE/xuiU6FPJLv/EImHNzwr4XRU8Itketj/uvj6S2tt+6NYvkPp78A2/sD
Q+Vynm+0z0oI2ZWWXncM1gTboUwM9uBZeaGzf7P2B/wno2DZF7RT6dY2eAvk3mdX
val1HWkUbIMn4TS+8JaPQCeS4qKUwNee7Q+n0BXw1Yqobtx0nxDpztZcCqB9XqWe
bwDSkscBqMUuFf9fYxFajaH74vS+WtIdg8uTB7wvrauifaoNltXbMwXNKNr/A80A
OVeVArSaELpcFMPHGQefSXM6SSK9lEiCDuox/2yoHMwiDLaCPLLOZ2W0EA+IxUrD
3yyNzO6alNqsEP8cHjKrwBM5AfJoJoXRLkCbigCtL6EA0tlMAG51VBA81tC/olvH
PcJSjK4ZYo/hPufYIVEkv1aueGgbCzYssBQAYMQCoVLOa+K+YHdetuNkwsyxTqAI
yr4NqHQT2I0KKstCZKH+6A24sPuEgXosAVnNMR7TlmTnuukkJeGD3WxjWqYAEgRb
LiHQSLrxns1NQUlG2ojgZrz6QwKQHTE7G7PVHbHYEovOVYoRJeg5WEB6DU/V0mve
XSKt94wofkxKwPkwKKxMWzYramJgrktAYVfHhbSfG/w7pr6g+/iJlMzNFWXdICC1
w/l16pdOTQGQyE+RKaNVUqLD98zyUUUeMp2BDJ6Lo9mbsKIEkNlwTPknblrjLHVL
ylhYsE7FBnVFXm/+H56fLC7FNYpssaWb8BpCP/nC/dptcFo5kQgOSaq7/qLsaAaL
+Ki3Ao3oFHTzoKCJ0CspB3zhrp2u6xYrVxfSX8xseXPsN1z3O7/uLcc/RvqPw+No
zZcP3dSIM8CuI9XPcjO6Tur8C8lWh33xpOTEKgO+0ipNz4AOYlZihGQAly1caRSj
DydUlJ9SisWK/cKeZDieFEc2Jsdq9OaRneBBbFQxYLWf8nzRjcwi8cnt+9UgC8UG
ek0IEZbS6F270ewsj0DO4CsfowNlRAwqL8u1j/GC3UAZMm7cN983IDJ39RCL9p75
7METuP1mvQMwO5Rn1E4Zho9MEh4IvgG7DxKKkGsXlaExdBqpjeSyhhuzVPVifzol
YS43UW57Rtsy9PcSccR4fakg96SyJw74tT5gwIhOFO9iZuSch4944CGhCvtWVk+s
tBNt+cTNp+KfuvA2WvMq84bTkwPHhlsF4ZbAADpJ0xiOkNQWoXZROWyBVYb+gJHk
u+DpITKiCOEkR4x9+X0usEd7va9rdggiqE9CAYriU+HNPZE9uvobXzWT+G+0GvQW
UlZBcm7ag++lG1rJ8LhqZpqyOt259X3BaWwOoP7nrWSXtiVivJUKp9YqyqPUNMC2
UKxq9arbp+cSh/N1OzOOUF8OatBvEnNzuvsQQWZEVT9j6pvUfRv7sEc00s5ERypS
BcRRcqH/Vy0oVZdgd9MDYN2vcHh3SBVc4xn5tgc/fwZAqAAUffVWyWlp8zcsIEez
mJi63nbSDQiDf3javxKJyoZDEQxldCk4JQhigleB63A1p1FcSqQ5op6RzjeOWuKU
x0hgTul2QswqHJiphPsSwF1vZU8MeRn8t03IZPQCn2lXT+xcwrQKy4WulvAd+h12
DKI9N9mqWXG3fLUlXTFfHBe7bLZFgSeNI6xOcMKDwXr4igYCRNpEHLDHNdd0vpFK
EkHrPZoIKS3d0z6vFXilwtm2PTIZDXulmqHD4BMKX4qEBU8Q5GvVKwejhMBgPnWc
UPpvaSsGy7bWh6HWdk5KfRyCJ4nKGQf9028qnQLpSld/cq4gohZVxVXV6o4Tantz
Rd5mZZlX//ENhfYkM80qtpCuW2B54t435VI+AXe1TN+Zrn8dVIsL79qMuR6EzIYO
Clve3RpNJikUgzVFICdK/5scFLroj3RHJAiXhs9oXIcfSLeKX/mZ/MkwtQonYd/A
juF0ILnzwOoy/CKH4a3ScZfq/m7PdRkp9V+SJFAKhaEeexBzM4zwrxfW6HXuH56s
TUfNicd9IZlrXY5IlfeT4Eg8TK6kCEBFmuN2js93wJA5a/Ph8cjgNlpgeNemSoE+
s4p0oTn5ItsiVQdwPa9Qt1uD0B5D6m9CsyQs2T7xieiMRWqvsLgQN03UOE155z7Y
8bhmjO0SSWtW3PAG2hwAhqvR4tsfckL0E8+hpaY2+M7TYOE8cO42C+OuTdkyX5zv
DYtiVWj8wMJlzFs66zmq37U4ODIGTUSZvBk/wmunqO8MB/q1u5C6bx69ACnWi7vv
Z6JeEyh4yoS0ibvA5MnMWu/flAUhJ3duH0Ygl0MCP29qNKO3FvMRrTQ2RClgAXks
wcXOcy/Lkl4wjcmyfYaJ+lTZat3PqP0JAyOLVee74qnL67BZq6W8DJlBM+OQQNd7
TH4CEI0uX9M8dM7Uw7DLFWEDz78BjRlOQzngS9KvamWCNIK0INhb17tu3PFPptjP
5W8q1qs+nkdUPWfILelJPEPeJzk0G9MmQ1dIHdTVhhUDPZD9hhUuaJM/cmkPcfq2
L8MTy1FPqOshEkmkC0B4R3E8eslL0dgMLNiz/J1Fi4/YdGC9ls463fOzgjv32hnt
wPAuVngLoNvqIhws/Ugxo/bndiEMIfApeZXsdrij9jEpugxSa74wRfn6+JtiRMoG
0q+c6VZpPbLwgglI1Y7JQatv5b6XeMzeX1gkMyinxF4xC2jZajfQuUTtNP3cvH1K
eFR//KRl3Ibyr8FpfQ/NJ3Q7ej1XShuhUrjBh0WFk6hIvK7T1g7RKSyouHTCB6B4
u61MlqEIfl9euQo5WmIiK3WqmVLhW72el+G4y6ePish51hLAXBiSn1S7KVufWdB6
xbn+WqOcRdeKhGPwaGADDXYTK4mDdne1Kb9rN+Nvjd5ivDV8FTsCQvDuVm3XCfR+
bPClqI0STUNcbjAY6ns5XS/o9I5FVZJ/Lk5O+H4b890EsQZXY5X0zu7eyW3UiD5E
/MW5I+KdSR2CERGPDO5q/HqnbfiLrN4yea6G1BiSZKtBUb6KKqtBLq+t8COoUjKm
I4u7tLYTQh4IsYyDz7bCxNCd5tZ7MLFbJgRh7kuJJzUgU6AukpU8qmXZR57qR4KA
/UT3SeqX5jlBDFhwYAkvizrR65hgdE0lfc0Hk1jwIKyfT5NkVDZoqWv60/pbDUxz
VC3OOPguau0Py8frUrUDEFuTtTP1vH2W+yRvM90HvdPBkHGoXjjOcz5cF/KMKo7l
LakdxAbfzFucEZ45ipcY3spgYgLWkx4yFgg1G3eyo2RlikwJHyAPQFRnmQ0A20e9
Z71n0Mip1cp2wFETlwSY1z+pf33RoZAxcdfGb+GbfzcluTTeRrkmvnwaiJtx7w2g
37roY5sJ0GHiP6IxoU0ORZNSyR04Z6JVyiIrBtrKbKJNyF8TpXlA/7q4Li2KY5uZ
c4Srmc4BiFwyadZfr0b6VIz43ecD00iHCoSt2fPIA9YRU3jhecsr+vYmrW3O3AT/
oPtoZ/ERcNiX3eLLXT4ZXgB3oBxMDHXo6qmlNwpXs5PtXoaFuZqQDKxM2j6jKozZ
ExHk0mUcOie4pKQ3GZWqU+z4e4KKTniJasVqxujXy2XkHhVCTe0+G/4U4789e1pr
ZnECkoN1LNkcC5qclYNDeAuoIslV3WyBVlAH7t2v1J5Yf1rpRc4jk7KVa4ahTkv+
oZCKOB1xpD+AmEJ+rvyI8C82xbxWt67wx0dU3AORPPRoBunq1gyFYFd22xBUDMYd
C/nW14MBvzjyZEOfdNK5IthAGSAi8r4avQwWkcvB2NfXpZaWcXrqIQhx/3UOHcQf
OR/BuDhsj3L408ZfX9UlfmxPlKYdFkU0G2N6gaXySiozYFxI17/pxXd8LdBQ/9xt
plHPXcSRx/OExltX2bOAkybuL4F/QKsOMbWAeyah0egLFPROTiYhBeWzUxEi95jA
1YS91yRniaV4qbGtvaLKIYiaIfVI65Tt9LGPfyh4OXQk/REXk8lOFRmYyNDMmPWO
Bc4Zw3rDfldDWkiows76Orq2B5s9IBLBhr8LsHR0ODXahC3g/vbiB8xlyzzIdIVP
EJa3VP4zbcwLalwNPjKaJjK5idF1B6+UsU9YOXwlk4Ew8SXq4FFI06AnoP5+ZQH2
nwoIUrgLhaXjyD0il94bkHa1xbXbY3UziaZySsrslPpOTdgF86+UEBWffJH24vnj
s+kGz2gksVeQC15LbAnzqmQX0Jm7tDYoJxtq1gc2JrFp8D16gxATlh0mEbEq28Ld
LlGGwIiRGWtW60KV2LS/HDiVdVc6xrqdZBPQsCXN/n/bB98B0+uPfU4I6rGyaoPG
yiuXLRj/m+iIYGKyzmGzTSgixPVr/zCRW5jRVgJYfwzdFfzZUV7/wde3gIXSteaw
VOv8nT7fayF9qhXxaWvm2vtj4TqaBFQIiNrhC2Olse1cAq93nrKGim4Q7wzEkQPo
dqJZOpIeWvShPhNRPyaQ/QhIKJQMTV3C2nsNbTDQPWB2qCmckd3cMaYdNNSD9hDY
1HDWC9w9F1HJrsn3U9+K4ZweSUNfbSbnOfqi4VCI4maNPDZEU/Z+RF/j/Ek68IdB
IDG9uF4iG4CjbvkBBMzpFkbitdTInsK+APgDOCnS6c11AqxVVcbGUH0G5Eqr/gwK
ha0obcu1wg0oIDaN84YjgPTWqX4JHBsxiAn4K8xGFyNQd4gCeOAIDrWfdq3I/aLi
7QFuIJ4Of4sfNb6y8aaDPwW8qLXZYuZFvubRS+IVAQSDgKoXvOMxdzPQjZnzq/Oh
szdJIM1OoB/pA+Md1lCuxNSAt8zbNHI4kfpGuzUaJBRah1rQ/98r2sfx1kScm6lp
xw34tPDtDfDdjA/b9i8av6Tj08FMN4TREBWR0xwiERKzDL5VYWpSQn4h1ZZt0P3o
AYppofkaxdsAT9UEbo7sxyp5oBTk4/TO8LSsjX1LzU8Vhk2BIe0kJmoq8Ry+E8Tq
09SKaWYN8hbPPf5EkOdgwKUMNDuQSmTPAixyWz1nWu4DpH4lKQRv/ZqusNGni7g/
2lk0HReVPvFKyG1xj4o1UhynZUHT0wqgjwOQDSzq0B5Ei0arYvVXCcipD9bw4NAk
28ASyVsK7gSuESIOCIz+i3D2DuFPP6T7dnPmS8t8J9R4/S+DW9MFfre0g2FJvgtD
5AfdmdTz5eLr558GY1HIsxU7phKQmeNjG0gLSfeXJ9/vYrpHA5glpqdCjJd4f5uQ
Nq+/pfeL+wlyavR5PPIRJxfgdRp+foQolT0N+FvtgrdgUr7jtqM4HgRS7htKA1jj
YVZtp19ipOt2GDHNFpYChlJFWVgOF1eQEyGsXD7xtCl0J53vf81Ux0VegXF2PNqO
hpcyl9t+AxofL3+//Con6e3otKD5xzczSJHdtVl7wgS2vRDxHpq6hnR74hM4vXNT
vmSHen6O8svO7J4uTsJxnTq4iI4WnxtO+yvZJobimwN6Yh+Hvist/dyEN7BPqFba
aL2LLsEteX7IMG7yvkKqTrYD/p9ylRWE9MPbd8USrMVsaRl4XaakNv5qP2lje/Ac
Sj43TqaelDAPzR0xo+rKRsudoiwJtNlepIRDbs9DngSgsuWt0uYSXhjbwPcjhFoS
eV67GTiDsbR0j+N19a5KT72ujgoBza1ii98FtjetWtSTt7GyltV9/DmPLMuf6Uq5
bn0mXrX1v0VNXxwnLuXNTSiCahUMP1/23F/htH8x9B8hVaP+sqp7UIxqAyv3yAUH
M6ECwXuMXK/3/C/f4YOLFNuz0LoTvV5NvLTnpDWn80UK7QRSiHzmjSOz7i7FJkom
ZuwhOfgeY1Y5OCMiTaz9uY6r4TQHS7dn0oZaRCiWVYjc2tm5akdJTWskEr9W3AQK
7siy3kFbXwx0alyPDA0CmrRlmHCSkA+e0X5fl9NlCeohpX7CMBhApzGyFtGVlWdS
0VJtdSrTtSmd53+JJ6bfY3qEaeU3bJ4xLv6jdzZGNiFD4t2CWy9a0gFMnSexwO/R
ZFh5AGyf1BCe1fD+Qr5+Y62CFa2j/BpVClRLvp5GHTH98zjNVUHx0+lo7cPInlNd
mP+HBaMNx+9e2Q+mbp1iseWbAntz5Zb+cFjHKjyMT83ffRQOwZAlYmoQ2ViD0yir
UK9G4tHLfMsBtmfG6UQmSPgJ6Or7huvI0z/cuS+TnxmtUhrYF8FAITuufqZ50pZ7
W5Oq6WrhZpsXR6THdJWYm75j6koT23Tbgfo2tsvcJFO6vVzsQdfQ4Xsr+Hepntax
pNFzY6+bIFmnz3oh6txDeagP/Gzqf9olW27ziaPyuXwpSqjbxlc+GbUKtJ8Fnw24
F2Xsq7D9ZFzqwDJ85aCar/D2NurdJOvVW5bYctqnxwvfOVSSBO0Zdv4WBuS17Eva
sJSqf0xGhl9fIdDmXchu88kOJM+zvd5LZb0wOQaOqqV80kZJ0V9SpvuGHwz4qiRc
WBZh3mDC+UxhK+I8x5SMd/llAjAudsztB37q3uZO777CMc3ktBXyvFL+9JMPhrRL
0lTUNQZumn6SAuc/qo1WvsG5wDqwMYh0SKDcGVVyFawjN2VyvaH3EOD9A8VnjClU
6j3yMw5nN1AhUqVep2pMyBO/YrORW8AaLV9ZlK5S2l0JEbomneNQidAHDCzHpZed
h4CBTLGxkJ1eU7ZlXM0gIRDr15dq92TR36uJCpA+4eG4rB2VPCEgScdXXRBfm+3I
c8fCtD38U8j6aHzCc+PEaF3w+TbCiBujoJfYkv3jdWEdrBjkZCoihM6yOU+gsK4B
gDg0+WyNaWmNz+mJx5rR+QiHwGqpp4QelkdriT2fW9ezAC6zm6/1e7iKp/y6V28L
fWevkuQ4kEqVT+2itvcsKEf1HcHfkA+JSCpesjO/66J8ldGZvNGqL5uJmbZ+dL9j
13rCDjZ/PGUbg684rWt+iGHjTz7Aw7ijUlmR4M0U8OFVdI0MuMKzR0BC9z7G+Nlw
p6m8/aQI+PxxgZUEM+6SIcIoPpyDpSkgxUW5cJEr45A0w0nW/BW6xeuECe/SL9GK
0zgu8qMCg7hrrIyCyWU0NeyPTjZMWLAmXObcyz7fcqF1C/YJ3bMfroAQgGPjdl9u
coNePKm1dKYDDQqi8UTnauoVqnErX4iIaTjRFdpVEjvhoHIVTS5nEgAJD5yGHwwZ
+Jmv9XWUB+ywDNvvgUK7M+PeJq4MMJStThs+rOqquTMaw5Zv0pX0bbrB0xc4haC4
xauQwfpomeldGflv56yFPOTXicDHuqipxdKMghVqXMX5zZ+QM3GCYtjG8Z7C6rXc
JjMMl7gVpLCzeR307/1Q9Geit6/AKrdt3WOUK9WQc1RL75R87koml07lKUqHekyb
u7Yg20lFEEc94fSSYF5ti7kw7guwLUtrjkoRZ5vSVSjDtpP04EwnZLDxguQO1x0B
H8pjZCH/5Rpax+0vytrTiJMuVBzJUliYTARH5beH55KmBt3V8dwH/Aigy9GwBZPp
1brFF16Sj0F4kLTEYgjgOIctayHiIyZsSe6i/juC214ptCUrGjChPKIZUu2FxCcf
42AMAlSrgtHqA2PABWoKb6BaFLWcyHXfF13FCHqIfVYX/NKgLLrVYjxAlqPyFZVU
1kmH/uxKPzAnqpIfJINpWVTp+nDHw9BPwkx5slb+GQLZSrfvjvp3isLbwZdhfgUH
dkzuvQHg5kAreOWsYW6C4nM8kQzUQXhcFc/KBF4VH6/1Yoy+dqqZRbUJiN2uK851
A8cjfxu/YnK39epTxIXUrYD2+/fPsE8d/Z+a8HyqvLAQswRHIlHe5c0iZyYmsIYI
5xnYwTqPc8jc6WHKohTopbXVmmf35zXaEly6g/41l9URjDsH1flU1pH32aDg7acX
DWc3UAbCDhfw4xAR1NWT5LQ2n/SIPsNxctmVs38T7tsRhAGyyWE/TpeOPZqnx90w
toPBhy1z40qypvH+pxL0sQoSUE6XHHu8bXaa0G8gjI7Gko6VjNb8PCvUIWJb1i3b
uWPVXq+Kw0aAEWjaqbvGdyzgFLr8iLiYBQdxngSy53wYJ/wYnMGJjtD5Qtf3AZTF
mLrw//P/YH5sWE4+/RRqQ1zdCGpEbY78oLu8hCueQBanhc4932OOIPSpQPcZBoSv
rvClNpRNSOSTpD/qL89k+G2NPcNxqEYmqvzyd2X2YHoT+wbJCjJhxO00STauctV8
BoeX2A6KXfT0tEyYa4YZ9/lOF/4rT6B9KHti3ugpR6Ii40wteO1mGZw2X9DS8hZc
bTTEubkIhDqQCgTYsY6pTdLT9IXe2zGXPPUUfvqG/o7vvktHngC2l7rm+dAu9qFQ
e207RSIG1WqY3I9mc2bOml9KAnQEqQEcvha9chs5z/rSslChOA9td4M4eoE30TzL
X47zNIDhHOE/KMgxv7ZuvCga5yfhiMRK8lojJ8tIFrwKoN6e/pfLLxEYz9P6lIWI
WoSt67cJ06EDajHnOo4y/763BV401HITDEH2vE/2AknAzWODMe9Pc6E0SpSvY4xf
pstKl2y3EaSUvWcF8ACOBaAqM40ABz9JwmVy0lcjmtD6lJPR4LM4hjfvqx4n1ABZ
qvchYAegA0hlw2CCKfGZM5GwrRzR9MrJ+PpSqRMRsuhtD5WrPlmK5vvTqn+RD03U
Bx43pKDPby2o84ZIQUC2ggmZ6Y7rZ3+ViPRi6TfORlGrdeVqoByArlvFaTU+UaJT
pFOtXDr46Bs8YAs0NAHHdWCHiC13GTWvYIPILC7lw/EY1bsdzFn0HPfuRqNXz+le
fFH6+I8lqUyJumjH9bE8w3bouTAPoLCjARkELGJ2HPtyjp+olt8QJWzYGgULxqpN
id/4n29lnhHrP9F1jpK24itjpvxDaAhM9ZBSfz3KjYhRZspKc6Jyk2NRMFLhp+Gi
awixbEd0NvrARvsVQiHxVjNBpmQoPH09QsSRJ1c4O9YyhnrDDY/aQyuu8S/tahJc
zZooA6SMoBZRfAtnOthC37mF63dwvbP9YI2I2l5pghwXogFjryzQTGiFuM0fb95j
xmIiKVdDudJ9eYY70q95IwZkte9L19KCFP9ZvTyuhqliltODReRAZH0WAS/VLFrA
ADL1mzy99FBRDUdZTe3aJf6r/4PH9cTOq3dTH+btfDmz3h/hWQUV5zNvWhM9XTMA
1WWHsh50v/EkiWrDDmGNcHDzJgwSj3QPE/SeABLfThTObKpQQUWWJnb+5uXsgKcj
JGlcsfVGTiiHdpQifrwHDkqM7HadVM+aLgBfLkbigSLFdDsHJ6eaiDpOnqLwjZBe
a0NPdMwQVdK1L91udITxqyW6Bfj+iYgFjJ71BwYjnSiSV0V8iruO6JcLPH4J+sR9
u417v9OlAAcwM5ecvoSy4CC+Ne+Uvyzub2RGeft+BzmNXsjUdiv0EWBrCoeQ60TV
qIicZH3SM1k1fQaaOF0qcOztnScfpW5TzEj69JWMkg2c83MEWM9oBLIVGdRSZZp6
JOPN2DZ6WfKEyECLHAEwHMbmZ027SYq239QK4UL221DIXAvaimBCMrnlosTI71oy
GJ221dBVCoEiiGA0viow5XKvOqb4YmHVBBqNGAqqGjjLMr4BvasH31wXLBuFQBmX
gqiOngKiuXO+whXgrw1knIYeViXyOUelgltmLmD3judoycY0/AHsaprQl51rOLXF
wQM3dzWErGUi3X3Bd2FpwIbD6vcZjhbMUrc58BmdVa1Iv+fQVmP+wxIMWHbMhar4
9FaxERvJdSIxkciAj7fA2MDynwFAFGEMuSt/WG3UnfZ5dxPGcclh7sugIOFwOibT
tIvZv9dISlUU/t76OoUpSd1uJETi9MBt4JU6JjKq+rKH7plKIDY2CR7othwXiFFA
gpNk3t4/STIU5EPxETzvzhHmw7Gcc0E7m+Ri38CoHH6KqkIy3XOiKk5NM7HJ24Rz
FJS52bdbpvOA3GZcuiAgCUOCpDCm2f4tgc1VzB92TNJo4RSiU/xKVnhnwejQEvDg
2mSvb+mdbPgAEg677cInKecmnpw2jouWcm2QEUge3QdLV0BtEK7jP8i/LBEbklkq
0/NK6m+hnUY1n4eU1jxqQ6408VZCZbBDksOWH6oWB2OQLs33EKJ29lAsH9VihbHP
3/RumlalWq9kqA1FMJLlWda56uvxRtHAa5NSlZc6XmSj8J0uyJBndrFlDqkrkSQI
V7dud+X7039CX+3vehxmWnNxcjtITh8fgm42xRdhtqpPwzvgNi4vFnH6MdOFom54
TYm0j31O66+w0mB8RhweadEXJWbDwMjEPLJ+Z1Y1zfZqND2I8FIhGyP3W3aVLp9l
N+Z7AcsOZ2m3vhJ7cEhRDfzlbD6LUMFyBT58L53YuwJvUrgasp1CkEGInjma3J4E
T5LvaIVqzIQL365W4V77Hc5+o+xiHv9Ki2iBD1feOaB/KApK8GCdB8TsXmSYGPIw
ei6LQsjzswKqX4/K0B+81I7hH7F/GEuvqQpWJ0Wb+/CMMdzVCDBX45DktJ7QtES5
IgroLanFrCFrIIfBQvR71yeuGBJ5z4oT/lmxc+9dnf2pX6gJU42HCsE7SsbPv+DV
UM0McvNsd8CFbah8cEu4JEDcM8X6c2VOvQAVG72/WJKkhv3y23uN3n6KJo1AtYOL
G+26qlUuon2hT+PhCIyJb2QPKzqAYUGLimqC4E69llqL1URdBidJ6m3/z7lyjttc
qwzsa5Qu+uAnUUY86/7NMPk3ZOIjewYSrr2PABeJBxn7O0QwJ0QQPT8i7KlacF7p
amEZvBvL+QEGyu/lru1PMV1E4IX5y9iI3kFNheJWC2dAOyRDLwGrsBN7DlsCO4oY
oFsgRo+Aotj5YjF4Oxv5D8Cl2mC14JLWAmo0MmnRSQe3DL+LIqR3LvxRP7mBb6+Z
rjsWDkMVx5mksYVwapCDr88lH2NE/fel5DQSerEVY8qj9B4OxgXQ5NM4GtkgmYiD
o5EJWq4EXBHzGgymHBjbB01vFoF6qpjiZy9urP3HVU6c7FkQY9x43ne6P/Euc3qq
D7nGt0wYhfz3a7k2Df5X9F3/99kKZjSNi+dPb1X4pZGcCEbyICDY8IJUnfugChl2
5lRZOyLcmAzwSei1+ywL/cJ7E/KvZoQ2N9px0tBOZMdquTT/WC4x4grj3j7e7RJM
IorTuMD4UIa23tZWRIMNqyw949wnWsdr0LOaa1EQakbspH9loPzAPg2ULSy+cfcI
lQZgdo6+b4aZEGAKAvI1inFO0kZVwA4JVtIvs+T8v3F+18rYCP1GAhlJRA3C+3Uj
Xo+33+KcicCpDhxLZ27Pd0xallil13L8GvGU5ESnjN9/cJp04USBILF/EpPoMbPR
U26yUZ4CESV121482j4J+gZSJS5M+7bm0ttF5OaHuchD9VQqHkMWpjdJy+DYoaq7
ZaOvdGKh0NSBLk9GYGGqPo3ZXbWwRPFuYr6RrQ4FKbxDrqpeLAomESBs4+dSVWJg
wAjiBJTqg6EED1lAod8b5v1sP7np7pJzfMeBijjbs+z8AZ1IqJ7juY/uvFx+9zWz
36s45BkElr0xWLtmDroQt+mc0VPwXZS7X0L2z1SwM4y+9wvBC4c06Rgq0MJFL8ft
oW1TD2UaODjjBiP78vBd7ydaonnlgNt6oXyO58Y3KPDrhIZPU7m6O3jbl1+k1Z5C
I/mi5qFUM+81FnIvaEMkeNuDZr8lXwsMZp8EbZfsFQt6IXEqXXm1Ay7owygVVSGT
+DAlsXYGlbvMrfylTCWEYSoeA3jgVzNQfIawo5CqYe/yBoEpzGsk2+in5lScLMb8
q4cJmOeNFRHoZ3uc1dR95/8OOJ/1y4QlTciWWcqLWaQ57nKh3MXBkbxg25IM2su+
hZlVZXI+keSncSqmn/XFoWGo8JOej5U0bwQMZ3siaOJPusaEYw2Gwrc/SL5erGke
yMtwOFqsB5ryv0RzCMXVhrH4mRRJwkM85v/Uh6TTngYf0miuH9bpqEKYtlgEH7+c
ZAJghJAVrZJZjXOzI7sISNeNnSkqYUfYs2pib8cU/MbYJ7xM64bAQlfqpIvHUmjb
iJBiE3hoEIe2ggBc4K1ojPOgBCCbtvCa5jlKZvNQl71YSmuNrsWikO77GspRFjVu
8ZDn+e0OdXi7JoQenmaxtuHcihzMrhyfw7cLd4RfLVaJf/k0Jbh0ttssoRFjsSsP
kGFM7Mgllj/yeKdY3s+99TtEhbPMK0LLCS1eiXAi3Sv9DqdyiNz+XCR3dswGw5FZ
DiORu02pC3uUrZTXBkb9DxuspO9rChOknTbBoU4XT33qHgr8NbQO36D6uKiiXLuS
mO6Y5Dr+B73uRbYSbALCnMpxpaCQj4EO5L/+y6QExuzbZGzY9ydR5tWralQE/M8G
R/Jj4XqoPbdztMjKN+5fdniR4NDU8eDp0OWUDmKJFfoAma/RHxfkNVqh1zxacPGT
rmadF2iWuA1v9mBJvfyEv2K2V/B79ORjRD7UaO2fcIXJKykK2sW92YmILDl6UiYf
EQj7Ab3Esu9UzqqxJNzvR8Hwp2AeUUfJuClPSkOPSqCRmKy0lkDgNkkWouj81oK3
pAYOB9QEA+D+QkDzJoaBlno9BdpGxcpMoj8aDayVxyYxe3QSihQwxwu/e/yQfiYM
aBY1CpK+0Lwwz4zeHaVwvnWTIxwgWQdTrii07OiJZywMIwhnjycK55Rv9un0m7He
2O5+GQxrYdewUcnnmMfhUfu9TLI9iHo8QIxuAzGF1RLTqpmJTZDRAguJIAEHGkRk
l8OIAXoQcXm5Bp2VjHqSDs3lILNKLJiWR3P1yHiHyPGTbopnxCZWelUH0mmIGviQ
Py7wK+AafyJzkMuLJYToZXa1w4KvrcnRP8IAiyzODArQIilJvOLDj9U1rfUXnzJV
4xC6lzcZBuJB+lDDCH4CgicmNPmAPqnB6+oo4UPRaoTKKadv5+JLyr8cqtBGxQxW
8hyNWkoj3+FsEmiZwb2KR4hfxIbrpchQZMy2G68nxoRw8sv8d5FiLSFD/Azo/JBs
u7yiKpVAmuCvXFO6R1XSdqm3VrRglGvJffP+rkb10a5TygeHVBCRzyOMo9J5SSJj
u87HnNUstxd8+T62+fWZ2cLAxL12yk7/Ji9ErqdPRXUNK1Qp6o8Ck5zP30Fg5tpU
12nsBIz76x4M4imVLzv0zZpGNpB4TfOQe/hvQUkGFRn8Jcn7u5MO3F9+izFf0WwT
bDehwXLGoPjE4F/HbIn7szUXDZMCfqszK5s+LCYildLDPxgczdMqq12kSjdhwFks
EUKZ9vvttAoPgl6cHAe2RVb9cS2HT7Myr7m3iDD9enrsbu9tPjcJCWFIoRMLn6SB
SVO1dvYB7yQ8rkb4pa+YYsvZnQErQvqMkr6UzTyKEsJjWRF3etEOrGWpazQ8LY/2
PDQdaJuN7o2j7AWMwFmhAW21fJiK8Z0Q8txl3UqKCvW/ewPjA/wjeTRNmzsSgwM3
+0VEyd0SdN48sJ9JiqxmwE0JTRW7NcZr3b7qkrhHx6Klr0U3SMJy9k7NKo/IlhyR
Y4JuqH9mjRcDZQhRLCyv4NN063Gw6CrN2H5fjE+q24kzWhwy8DNc8jau7xkFp1lu
wZK1JJXOHNBTYxX3eWAjeywr1aSJ+JMgs/DGB495yBI5gBXdDvB0LZCg9VMstXZp
rpKpykCl7izx7Di+6orvwoxWtOg1pr2Tbm9hlrhj2+DsL11xSMSXb+soUpg5JCfr
XZY726UG/KhB7qufcVVfXBdELFWGvwlaWj6iz3bDnMNG66UID4JrA8wJbY+sXooO
Vu3ttioLjYu8uu2Hf7bn+loCUAJmLh6LtHo5kl3GwSCDSSwJbbGxP6pF5Vo8XOVq
LGnGyogdB63DT5ZcWV7B+oNYE9WnpSwl7VdDp5uewfgnzyDCNzgNiBou38/ccs1Q
fm0EMEz688+R4rGg3Z7mYIdfMg+3Al1ljLFtcuOtOkYEGgjb/tXHh1Q4S9uaTD9j
1qng68lMBo14tHZDIJoMuNTMeK6/NHGckcNdmGec+FtaHxghKLD+HKPoJ9gIhsy8
9QR7Clqvd0/m2FhRYXIrhS7ZytBw8YHWizyS6MuAuy9+v8WuqDZHwiQUkcLK25DG
hnT0mnSO2Lfc4aNzkpzD6MqnJg/Tf1Y86ZbX3jHXIE6EC6fABMxTR6xk4Qd8tIvJ
xgKQOyk6w1o85lUABUnRj26kWuWjxTHQh+96hhlymglYmn3O+0kb/9uTXp2+VPQ7
vP/1wWRz74n0w3Pk1BQUbj9d92zi6eeODpUfcnGZ7thbYNPNCBfdOoOkKI2BL/md
iqbsUt38WXq/wGBh3difBT4zUhpJlT9yMRBMAk0OjFXSXw5LhU31YO+czOxjwzF5
/DiCVjGENkSCvkkVcn93PXHKzuB33CQ6Kijx3OW5FkzMDgjuJQSBjApYFT6JRutF
LhDE8egJfm9p83ONF78ekqMwSaJA2wvdAqVet/M7raFnHXK5OVZhVVm8mbZJyK3W
fQOXpYHIb67wAhtyjs3BHvsxsEO/IuvebC+cbAGRJUYxPgKKusVrpBOBXB9hLdo/
mXKc2NGPj1eApdL+rP+gzycfSebJ18D3oCFE0OEXPZz5TFASEpVqeVbGbTYNLnUC
VvvdBL1ICthdbR7aNJMGxSRN5d214yRHW6YKBxOu+l75V0LmcY00PkuZVa5epRDI
m/1xV2qr8fsgUlvM3Vi+bUk5XoWhlYMgJ41N1p96YcxvjEdNk6NvoU0vD/K//15q
sI8fGLFc6buS9JCIOEuclCAHfLE2AOz5JCTfvmCQZhhX6yPIoI+K+Bu0ikHw01vK
57e4KuEs1oMpzfQw790ZpvmjYwrL0XNeQRossWCO/jYXzI4/LzrrS6oncipjV0mP
961c8MUsYVmm2c1IkwWgeMhlFz69Noj4kN46Ey+9WGmw4LGzulYwdcZxCsyIt4U1
VnFtLZleWfGfSHKyPXKdjSG+68bOC5/NgmPHhdrt0x00u9jnk0/zcCQd05dx6jdm
QOcUt2ajw1RJk5mnJyj8fyew2HB1Q1i4+PRWf1UpOTvyGij16RUCd5zTbPWmlV3B
ABpt8cwGAxoFVvyyONgSs/lDxvrIRQ8GfUTc6O/DFdELnipAMrsyJj7H4eRYO5UD
RvzK3yMM6DgN3ikmhneubZw5BNveuVriLB8MH+jtbT6G76p2GAtzwHFAiTdEqTAE
SpZ3CqX/yJNdFypM80jLN7ndSmZ0r9O0UWJwW80P5Dp4aCD8/kaIDU0D4eWveo7p
NtGZtuzJceRXTovj5DJexvpQSwQmQHiTXBKZjSpdF6E/8uwm9rtdlELPuddypiLY
7zJSBTns9xJ3HPy9S+khKKWtIG4EJWqN3h6qoPku30VSKOYVmoT6igtB5nKRwJy9
kgF44hbw69t1YdpmFzbq/BiBYprZqq4afvI6AL5ECOi4REmqRXICH1anie1dZqui
ujqEakEz/whqwYSd3rILJ8O32du1AFNuTPWxq5j7TZ1jCiOYYx7AqdvRCSa4YmX4
/cHNg5AfLzD65xh2pyJbZXVvTmH3rcLA8FEhcFvYX1+C/88y1joxptq1IDffLTpU
Ggovx1SsRR+iX1ibyuRsrd/qAhwo6yXiQbyg7jMr8/20QoESbTxMB8ow+czmcGZt
viuPhSM0FtX3XR7FKlbCSc8MkUi3WHbnGL7qYynXmWefgWIwubm3c1L6NE4I5CaR
wSwCC0ER7day+IUoGXJzj2wt7hN2F9mpnYuGu/+JELKf3ou73rgIygMYVkzJf6m0
/GYo7CeGQ93ohPUzFi+maVZ9yDW+qy3tRg7L+jVvZ70cCeXz06raZ7PeVaV86y5D
wkMT94q5SseXuyz7BA3o0aotClmY17kELM0S5kTI7C/OnTXt29XoCN10QkLswGod
IXn+RIgDlsWQupckT6TqNQs5pyVGwoKs10YQRqtW7AiU41FzFCGL3DFTwzG9IjA8
Lx6Yq9ZDr5lkPp0QHUul30oqeC/NpupStfCu1Y8EFRBzsR1O6efBpxJ9V9NhNTAj
/F5SItbzi1p4hLIiB5Bcsf1idDCAyuzJ0ulKQCYVnjl9GE1beGbkSPwdYtPztuLY
EumsYwRmXf+6f0jrVpQ7VLIxxaL3AzW6WnmBH5eTLPXgBX/VQv60A3LdezKfG8my
DeLsohLiEebooSCirowDuIdITjfg3L7Sbo91+7XkEbT3RpN7iO/u9OrxQqJJbMhP
1hieywMk/jjp1RYTQJO8WQKeRinclwZ/8OuoZWyBwKyCY0SSDuIo37Q+o6DJ1tHv
iqVIwddPrI5InEP46DrW3QVTr+XKiyzrWj1PRGJHB/gXjDrc63eBliF6vNevwfVU
MNHPOreghbMWdPa35g7bVusnO+nmB/t0CQ4iXy8aLyoGZSm3VMunVkya7cU8LFg+
74u5iT8pp824CUygnaOvIDZsOPbcjundStbm5wyHcacW8uMeZrck1Kn+yFLBfYel
c9eTOQ5fhq3sxIG9mxUJKBseB15gzCA12XTMEynR/TD8JTliWC0XbbKRjM1tYuxK
JtodU51wKWxDzG/wrH9KAgXQxRY1Q9WUU5Vy8jSvfYtZjUjrIGAaj82l8suN+FQl
tMaLMTT2uLoJEnLs1/IZ27ImrSQKMqTWBFro02VqmN0Y0L+qrb8DlzXB3Bs7fZak
OcroySjGtyBGAUKldjSv0SbBvwwRBfL6hPYl3T06VQ0DAA3Uey9fRnVrqlnqhXSO
rianYPqwEZH1mzJhU1P/DTTbTL02ljrWmJeHfSqFqqrkaADkAj83APBnmNmrpcdz
5CX/PMHYofRo7EHGBfzPyiB2oCOfJNB4Vilzp4IjP8dKqRQJNDQhkyMOm74NGn5A
/6mebCf1RS+aORT+J1QKjtEH7DF+la5clDa3E866chZxQPxPHynvMrJ8ByHBBJYM
JylXI21Xb2WpcSn/cwnpEaLWra5ZCBXG0hgZbR6JGUoSgEoX7gmd1QRLt2s5wBy0
sIKXxVDrYbfI3lskj5teeFFDleSmDmZMqompIsA8yrwX8aZbTPhFJFXhArXsEAVe
j60U4lZHyLrNDmXx1DPSQRV3csa3Gk3QIgLrW/K+puidaRdv0jnRcIOojvS92soc
3hcg9B8jfRYAPpazEKbZZS2Hf5/rLMGJiedzCZHHIgTuPeB5sl0ygET0yJUSZP8h
CzV63Y+oH+38ET2mBJdxOUcTdCFchFeSlYOZPSSC4iGkyPjYYfQbxtnN3bsaTD9C
sKEwx2ZwhyjtqkClScenpUt7LHbv3liY4CHAEeAH4hf9ckscQ7lsk/rQ6kiuoMFF
biTTerDsB76I5Y5gRhSQ7snqF8C7qYik5zuDLQhf2kZJ31U4WUToivoUQ/EnPLdp
xf17Ac65GGgGuk6jf9s/prtgwTG70J2UdQnhWIGsbxRRoPnFrE+7fcM9kGqDdgw1
Ex4pYmBjjaFNb1u9nsVTrmS+kYMnmaqJZfu/NBn9MbO+xcXAiVZ4sjT6wVTAtGGs
nGDDCfM5Fmx979u26Y5NC419q0YOw6EyZChSetlwsH7PT23MKOg7uO8k/PnR0peQ
gNJ5lgDBZfcXHslwsYAlG13BFIkKKBg1u657YgNoQmwVjWxr1u060pYOM0Hynjzf
uAkPJTgYPaY3iJa3rPSJwlBqksD0u7FsiUKdlgKePUEogYD4P8EP0xsYaHP3EvF/
aXGdJhJfky5VsrxjM4zbKhbz5rHnj2fCBWNqprHoyxEdGjWQkV5ojQp4vY9EGQW1
ydqevxAihVQKHkNKUuEbdisiwqdv4x93iv1zuhXp+jWgonU5JGcDsyuF9I0+c2L7
7rwLwhWSFZ/+JTziqbge+xGbfA1IUTSW/BVuABQ0nhjXcWnZjrffTI1PUH87DZZ1
Z0r7TaKGQ+k4QV1exDFxnGeT2dGHnJe4RtT03vmPzZXSPO893VVkdK9vChxJfkuc
eYbrejrDMst4ipHiyg9xYMQMYywiricRe5Res0PMk+Eww/mwRcsGMrdVOgefppb0
Acn75FfUco0jUF3QQiqPwju4p/vh00/MnHF6xyXN9MzPn/MWdRLoHrmitnn53kVu
OAFMTlRRjwpS4Kd6pyoEaFf4ekSwruJu9SSznGLnNDBwnybmMj11axC5gaAqaj3E
5Jt8JcsFmp+8ZR+vCpRB/pX1fD025DVv8zRmuVOJuLSuvwBJZCFRn2f0NG1zuC9v
D8VemkEPxj1Fkn+o1qAIIEvDR63hmtc2FakQxC764lbyzDsNgwncpQ9inTiSzSP0
pMz9j8i9Wp2EXJ8NfFchwuYVRiGsMb+y0ciyEinCiFg3QdoZtfGufkINrxTimVVv
skRjejZfKdXdysj60suiBY7aAjWbSCjQ/T7bpLdZL6Wtz3DX2oDCEtTZ9cSl4RZg
kjERRpFsS4oYqTUsNj8OvMGV5C6yJ0sEWBr3gZxMatXBGQ/BU8+hHTFOR3dh6cVz
BuLeDiyI8wPYjmnsbzdZ3u6F8AUlWpcLBlpMrnyx6VkCTyPjk7WCXtqw65THa1SU
wBZWDoP4SaEliPhozM33N+Vc1HmDAqd6v/7DePIM/W9mTy1m3fFU+kojzINVEf8C
B0NANWmKfF2AfTDEFWuJajdQrUqhyl0Cl2Kj8MVq+YOCOByOu048sJyFdrxQR+uH
If6MAB5d6OgeuKGPnNbGAVgOFuOZhlSxi/KCDkMyewsED6gTpHjdHNKcOILcgYvq
jafwP7KiRQ7TKteODuK0GVPnzPBJLGKuCqPtE+0meiHx8e0Nf+Wxiog8EE9AEJy3
OBq2G/sU2zqZUPtuO4tHtz5FwzNzPLwf+dOsCbRHx695Bd8cGQ0l6iB7W42FrLAC
JshxuqtbxP5PClF0UbkrcFoTcq4oXvDbQmN6NBR8+Lh5wd6qhRh5c7i7D4ztxb7S
4WuiaSWhcrr7x4cXEhtj91aFFkmMshdER41Ymm9fm1u0+tt6yO0vJNbfhXFoYEvP
u4ZpomWf6YtGK4zg44q06UyEe7AC2u8UNv/td5yL9iJdGQ+Hq1GWzsF+m/Jpqtzg
8bX5v2BKNC3/lRb1V8kgsWXG17oyOyKM88SWk4blDfV2GxBtUzcyKheb7O1ePyAo
fIu3u/SpXulJ3jaXFB7SjPnNb6d/Z8MI4R9ObbJ71/dHlPv7Spd0GuZXbkCx2pR1
T4WFesh7f5svSZKxDthH5gURifD4XwlzEJIti3vId1PSAhu7LIfJ04fPh0E/PFUQ
X2yLqWiffxngobXcVqSG321nKppvsic+syP4subfDV5qlQ9i1T86o1vxfPJzYRfD
SEfV4pm89p3SLzrmHVqIPY+/gLmeD1FXhvsgzXJHcBIU0Lw08yEVrmUKBtDj9rah
E29p5JVWxIgYc75oDBkrM4XXTe458K57O8su128YtxRPGT3gq7u0zCBI+n2LgMwc
nY2haE1Ymo5xhY98xKpzJUdQ8WnEL/v+4EzKS9X1y10Oy6N/xywxTQOe6n+XBTp/
pSJ2L2JjK0nVhDGb6doiNajD6uPLjcsk5CwCLciTnI7IbpLQxI9dFQDFO2h0zsS6
RorMcqK4cDqRF37dMEX/Mxypimo2ErPWfN86Jcx6EpndxvidoaEL4UiXtxlGdjrM
nYspBSW2nV3fB5ZbY+lEdqmoYMQ89cicM/P3ApzYLG8VRXyq1Hxn66Z/dOLPw4hF
Bi3Sy4iaCdfD2q87/h4thy+7NAqBWVmRaiiS0xm6PJcOfgHRI3OWK84NLz+Y/SdM
UGG6nqzjIGxE7DBJ/adnczHtnHs+q7i3u2uzZPxexx5R5ekQewbKujvQLYHXWELz
dTWf3LKrRZU/XItscejHXlE39MD4zCXgDZnnENRdFo7FIy30JPtmK0zp9w2s6ahB
VB4AjeoPmpoQxOU+X7g2mqOVG9Nz5VLIHvnwpd1c0WtiYlV9bFATX5vFSPjGfTVu
LTVze3p8owgrdnFseUhljWKK1v0sWI/oKqBssQo54LHKPwBUm6J1bto1KXMWXGJt
Yb0G1gTIOsY6rx3lMZbI6cVItczDVFt1o3jQSFXeX+dVcr3fpS5Eg94Yuj2/FIyT
V/7rzr0N4d7eLGyeuvUdLoUVMBIySK9OkWXu76Ck6wKEi6QSQ6l+wcXyE2F69+ia
cZHDRL/41ZeUahW9XCEbbeqDBOWMLDY4DLy91Qz9+6SQxnqhbm11hmF1MkGlBADy
IjbEqMLD83eJfQJllMtmWIpCuTk8mhyFnAb9EVw+DFEjt16ZCC7H7zLmn7XIS520
LmrLnzNWMOUV9uNjmS0bzRrrToCD5NdNq0YFhwLoaiQMJh7ChZYqx1/jZdwhmJ/i
2EBHn59PHrWgJCrk8eRG17PVi37/Tl/ZrBLbqeijMfogq9p8FxB2tkWrWBaXsdD/
+wPnZ22LKslh8DPMCpmKoT2tXK2zg6o1tD22BdryxhGVfI3PQ8kZZVQ3DJE9fS0u
2YsG4+ICun66NeUMfnlUPa0xbfA+r2+n/5WqLcOoOgwTacvzvIZHCEPpblMMvbKk
MScLhJfGgUQWwy9A1DEk0/oyvYypHvpK8JjDRESv5zctUF5tYuq0PiDGpbibky9n
IHeIonBc9/EgB9OspwQBlyB+sW/y4JLHi6j9yEfQ8CMhWBZ3oQNPa8oigo6BKWiV
aB52QWvrWBWKQY/uyjV8ImiRxb7+QCnJi2AUjeB3KBwLRVZCBny030ruGqnABYXp
54fOpj3a6nPCqkWOlZYR5ygE/Fl94V2unf+LvjTuJkUAvzEDz3b6UU18jtpxDXQ2
o+0rO6b+IovozY5MnT1Fchx+anzk+X42lO+Mk2kHoXVZJGlt8Y1a3fAQxZLtUVY9
vFbg1pZKUZ/gZnu2uxDcq6niHCP4CWYZEFthHDz1hoyRNjHuUvZO4D8J46K/E3jA
HppyP6XjoKw8x/big/Xy2pyZEyLZJ30rspWuyFxGypEZUEmCeAtEJSFTCHhD9Rh8
Zi5LbIOVTbqKhN428MZMkHS3t/lAR1pgB6+JoohjLespXOItRyHqIPRFCXZ+o5DK
ikaCdnGT14/PBppWJkL6rKXWieEW3A/U93mfG8NsxTheRSToVt/3mi0baJc6bC2w
B1G9x2IwIzuuNiQrs+xMBeLJc7ISQn6tsjvZRICO66K7u2uVeFx/Ev950fPT4wKf
K+L9DIdq1nhB9tjdUWruHEsxlE2EGfUI81XHc+phYmM/JtQNvUGieXmxmqx4vhBx
USamQGXAOAG8VeSzJvPtdcb9jpdj1gFBvxJWSdLmiwmkX3Tw+dRB6QWMPG7epoe1
XOk/xN2vEPUNWFjZdpTUUi7KqY6+L3nygE6V1/lKcnCt+xrl56AvrUX2Ivp1jFOQ
jznJZ1Z1opyzr1ycGnxSUpMeeCRjUYsI72hMrmx6gWYnEzCJbzR+dX7XwvAkxRGq
HkpHE//EWps3TGUnArQPsegYL3QAp7apc2JUAgQLdF7+gVPqQfyM2xcqXrolk5Si
jvmTNLBBsIGACfI+9wp53yAFW3Ha+ifNmprZiFS7oUKj5g3IKDgSWtLDTrhY4Ok3
Y7uotmQ/xNIj58qg0Zezn1l9ITv6Zb8S31bm+9A+C3dGmxCsVJof5/X0zA9uYGUf
IWhZcmulOALSXsvTd1cddiEXBNnQWC9CbDZ+ZqbZIVtd2i3bHBK2R42uu3jl4das
D6EplLin+7QxiRd/iYoI96rJjswOTjkPSp32pbZb7OMoL99UtynMsvKfaD/CKExt
DAR/zSMZKKQx+BZTkcJoze1v9d4o/fV+b+chIqjhTo5yGhP3FDrNHdNMuEPiC2aO
N3UiDmy/MlNI5T4n1gdt9p4lDc4XKfjlMR4t1RvG27072jyyl4joe/AEVKJzm1OO
9qUqAJg9Zv0lVeETjz6iSj/cZkE4Zp5JS+cgvRMGQYAan/0PUQlufUqy3ovMu4qo
K0cxbux8UNY3BwmXxJ9FHmGSDR+ZkWx9vHf1Ca1rfIiEdWSStLqkc+dlAhYq5uf/
VlZYfEvIGyQFO+jBJ9IZFpmzJW40svApBsQgL272DXfCiPrEwvfDKYzIyjD7CpIk
Wk8032tRH5rCXYErLFJruLoeoA0FdANyQTh+38zhrra1rtaKOy4nHB2oaKQ2vJtJ
xgG3G5niv47YgjTRWZh4PBpjGgi0OBg198R9y01/UXdYkHiyovJYeR9SW3yXQ40i
tNsae7kkW29gMF4sIzgH0+w3bRB7umcLKUOzAuYv28sS1wxMHC+CsCX6FNfXG5Vr
43O870w5Tho4N1sEff3q76h4uDV1XwyM6nK9vx1RpONZuYAl4sEo6Z8QM7Z+P0cB
5LY+BZoaVZHGlw2eye4aeB8s9zv3WZHcBYPTpk1KfzERyY+c0xbOJIia3FY1uLEH
fDXUGGdNHcxGtfFqHDdAY9xi4loRw7b5cBU8bAJzoS9Y8znsfmE526OQp/8y6ekV
pA3iGjtTWZjYVE91fGqWJKoEsfuUTkXnBZFC4sWBLF026ROEC+fk3VxMHVwWCEDd
VopssZioex0gOcKV6kcSAq/Nm86tfAzn0JxF0cNB9rfD3b9x0v1U9y84FQ0IfSWz
wP9ffrr4XHf6qI9HtEOQXhC2Uf1FFavCCuKajqt6BaI54mvFt5BGN8fEbPXtvkFI
hwhMRrs7r/LDLjiiHQW4jsULv7SvXSqg15jCClz5RB2rQFuggiH6aOvNlthEzRAS
zR2Laj3v18g+IM7nMhCKY8Ex87vXFzBg+cLJt1P7J9inLxZEsAA8w9y6TOqy6Uhh
2CtVCij0/n97q/FyfdBQADzztqAQ5nU6BrvvOD+gwWcCKUiaIvd6ONZHh86iWnPD
UQC+2I+DOKAh+XvyyM7kqsZopnFKj3WznzoejB3keK48rvQNMO7ouoy5a6IgnHhc
pzwg9LuHs/LirZ3801Z9k2EC7rY/ZYfm67//55oSQcb+CFBmVd17G8dY+YPWyUHB
Z/+ol06BmDt76YUF6t8ZrHakoALjXEwJUFysj89XMDH67TH9e9HMvuFqnEJ/TURe
dJ8Z/yYHPSGjlzP8nUiWqZ+MwViwCJX+dHHselXbTg0kL2QD0GBt3m4N2h9ventA
+mowpik2K8XYb2OKQ3eqG4DNjUzP82kOePtK79lX9UNscp7iy0E0ov60K/pHWN5h
bNd9AZE5lqS1prQHSaa6PBdYaCz7PYEsXHrk1jOtCup+zZS67ugCzvvCZ3QA1BMD
xI94CFX4tX/PqzajlMW4ADeU7KNEVHavCbOk3BPFkGOVsxzyW6B+EkL+tX0XxrOx
vQPxcy74sP0YTn73PfUJEaCfO597QUiZc4I9lC4ftZRdqsORjp7PqN2YrnDL+Hlc
aC73eVA4Q/3pG79QXXK7rUA+5MFTKHLxU/147S9vY3qVo/PvVuE5SCnowbjgvMZs
X6axd8UhPWA1BH6eBwO4F46ykNOZXpsqT8DQjtIaNXChwIyI/iKLrulHT803VvoT
QXYVtiOA1tEZUVX5jiNrk9VCfFxKoNNrdxuQl8lszhAy3acBGxaUbI10FrzeDaxd
R/9LTUPHWZVZtIr4z1+Obo5iJNaRtpUA+PaQeH3Wh+O2qIEammeP9MQRFFSJmSmh
vIG8k3KXq53CW6g/LsEIizR/F+blVc56rxE90sjeF/pzLF4VX7gVUfg5dN2hB378
kZMM6QvcOVaJDWHTFKS8hDbr7AIqj4iXijP0Y5SL29sKH/Sq0vxWH+m8E34w5d/R
DKPsLA1qnrefA0Xd2y1zkpg4bRaGX+I6f5U5Sj873BeAfROwUYkIPmjLpOEfbHO6
vXcGvDu/0EzEoGgXzov9VibtED8o6TpUkyQx4tSJdrQbh/JfKhraltfqs5zuuY9L
PjEzdb/CJr+t3sVa/ygJpnVsvjFHJhhPggloCWJbKarsYB0m+Igazum6sXd+atoR
+FTLYxvpYsxKBTjHMDuMUoC1f4CkkOBxPjdaLDTFO85nolsRnIZt4ZrvR7x/Vg97
HiR6nC3p43+wp25GNKQ+htzCuvNsx6QG2JMF6qJ/h9BbHkinvPOj9BQWnSW+cwoL
jpuOjbYZ79eyzu7bmxys0SGJMuGA6OOUeY2lhfPsGSm5QboWwab1BNl2msrXQs8a
b2Y48oIy7A1zYF6ZzaBsMYgHW7EWvVupoxHHrkwLPONvvCkWMPA9Y1ZQzfJct9hz
63kcpTt6BH5CTl2bQ3KCtWqtcfSmegj9Zwx5O76Yy9trHjMbV64XSdD43j0h1v1q
JYZm3jhkuZnkPVDZedS5aSx9l6k5quRb2S3ko98lJACMF0vA/2JVd8BeLV6htxfH
7HxLEM7yRQG2s8HJ2zDwb9e+KktOjSSbO8u11XYnVnYrcGcxDKO7GoQeo44Gn+ki
LOpUk8SnQc8WXBMgpbQM+5c15TXDKAD7zZxvUlqomJJxuvQKOmIexuob0byVfjkz
5owKAvi+BjYXjb1umVYthEjgM9oJQ0au5d91aXqIbhdXj9OFUw/KrAsbEgbBGdLL
oiAfvo5exkBIdBIWbAZ1A/LeEzDAsieq6pACzl4H3m41qvtYol6o1fMyMALVNipG
l/Dgr0gm3ESCicqP5AwroKOsS/k16Jo1/SnlbApXvENpQSDIATc5asjpfpMgyJAJ
Cg2FDjvMb1k1JkxhiJOQ1oPalabsXwQAGQCQyi5i4z6s7HjfQGow6i/J1JyS58qS
otHlg2k+0YsWXb3BKSYHuiPWt8iom2inDeAM7hVGUWPPKGYF5biLC8j6g1DivKDU
v6JGNRuXQIToRou/fY0f+DA9jmLFFANod6MHPZmT2J+lEkkTuMjoHlEgU45y8wbr
ebDcW7dyMHTkfX5DGkw2dR5j1fLs0dxJJ1txUDH1VYcVdLc5belMSdmME9JE8DyZ
UcorjGeC61ho+8KinyEfAYsUM8fztIdgSZwY3y/ezGAk7SQ4VNFEj2Yjk/zleUax
RYMylLjF5Sr4yPaGxP/QfxSZnPOWvBUqNHPawEYAvtj2LvZSIQylYBV/6uYjo1/t
cUL895B3IlELFCI27XTMpB/lrHNrmr9L6fVE+TDtjpOVt9AU2T2dMJveDYDIFbTq
pofu4e/BljApuSAj2MKqE73EdBhAWSS43bQwRotOobb6AaVBid/7HO/zJhyuSYNm
YMb9l+3HyiRTH/6QKFyh2qs29ZuCHcpLscW8xiu86HLNLxArWUQecfK2YamncbY0
a7fM2PhvAOdtaB8uE0OKJWP/sCYVXeobmXD/7AXi+kF9nVREYtS1ZocFFo93SSjM
YjYHjIz4d97pb6GbAu093SgFG5QpWA8WxaCqHo+cMSwEiMAATuZFGOyTwugle3yQ
BNmFJApEVEnTMn0zFEFA2C81/Q7xm28nONSM1/SfwtQ8HRY5YXA+AT8IPtZ4vJCq
XcENhgk57DWbXAKSvnTn1+sfHrnr+7Ji0+MMOpZFRIQtx9bzY+/FrQPEaTX/3ZII
lvnmN3QdYojliqYUdP6dbuzn/SfeR+FhPTVPq4yFVEv/UKzcMpVciQ45KWjgdsuc
2EwaQZ4lp5gS7eO//9CsAa8DPzMFXM1pI48SNCXUyqkWft0TsgCda82SCybSehqw
vtXbdLNBOiMbvb7j1x2AcMUwqeqn46RxeAM2yfxqKo+reaV17Wn7bZTUATYDc1Lp
aKWbGBdsZ6+ZFun9ONQauimOg8RAU9NW/AgwYAiPSX7s+TBUcRd4GvFDtwr8CmmC
76QEN4VCvoqpwO02P9YC4pOd0NAnGfZmp+Ce8NleZb/0Hk4/+Bt0MdYdWud/faqD
Ja65P0qrG3Xp1fauX7z11ZBKD+YpUmKtT2bRtEaCRF2Wlq9XrVqUTbpKTBzWXNpZ
lgEKpM8vK4iPKplVLQUfYYixGiBvLKpSZHguVVIIOTVy93zBJYYWF8zm1hHCyG26
VT8Its+MPcnT0CpmuXtdJl5SVHejYL1YddztXJzdujxl1sbp45AkJKyCzzAfvVHa
Rc0ClHnLjvyrpqNQtaQwMnQ/1hRaXBM1qXff/to6MPek6m0UQthSqEUXTYNyXNNw
H9cZJreOlyFJSBCWfXQjgY5VEk55cJvOGzzW8mxun+EdY/ibYvMo8k2pCT2ywHGz
NUJVWReyH3d5oLg8oODMU8rQLBT4/ylWZOsnsxwsIco/SezI4+XcavWnDC3IYNui
kE3yfoCn08frzz9tPKBubIaS3fHoLL2A0gwRdmP422wt1MfcD4pE+6oOzx1L000f
2CdlGZoUtVifFzOnAt/1WF4fYuYeJ1/DlXR8ekX1KaM5WbwW9tqIiaPxEgxO/zCN
q0CAQ0IYN6WLSVCis4K+3mhTf3EnfZqip5d+FcFhkP5l7ZelFNgsuUX7pzsgV6JT
Tpwaitr9Y48oetqJ2s8sZUQtUCo+6qJhWptAtUovUPnQOHqQI0PCr58JYs6z51W3
uUX2G6SPDD+Qwp01HLI66MptFjApPgzJu+m8zicyUKAM8FWpXMKqXlDBIM/V/6Y+
t4G4ShNYeJ/9vb4SXgLGSxjM28alC9a9yd2F0kAdUKoh4hQSUFEcM1SR9X3ddTOT
edIbxd3YEVHw7nel3/gVS1EMr5wecObQKsjeRbAJU/1xOpXnjxC97tXw7estftv0
OiJ23ND6E8bnSL7MKlWa0KlE8VjrH237CY0zt/NLvyVM5vOo5sJPu4ffOJA4yiBi
5Q/7jr0QnH1YolP19zjrQg==
`pragma protect end_protected
