// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:06 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
euAnUaV8Teo6+MKfVMe6lS9mzpfOZ6g09P/9cZcwwJjGm2Xf65+0myEGvmoueYVS
uB/08muGl6kZL8FTMWL6o+gFfAxMLB++1XEbvLp+J63/sIZg79xj7+DJmxnVP9kp
2Q/FhMhjWzDye5x/+qvJlwId+WA2s7FgL798hzQXRn8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32784)
04R7Agt2UEa+L+Hsamh0TbwZgQ+qTMYIW5H76pvwBCtLPft2faKeQV+kU5DIU/Gf
1O+2940eTgNl+DGaQvraOrDYLqFyyr/2b8S457u6auxRovGWM26I/V42UfQ1Gbjh
Ds71MaULaZBbBxRzRfMx1AAMOtCPBSbGoGmV4XpQVDiRjSO+uEdMaKQPl7T6YBGF
IubxKJDG3QDh2G+mdUCiG7MzwiwdM2w5oZJ9Q+h6oHRn2DwQIvJrCzW8w4CxcVVo
O4MmNB2C0YN60flYz+6ek1IX2uT7wWJSj7jlm5C+SBv1lXTZuVvooaaDUIUbH+de
OKjwehapHxwfJtZvo2nOA7IIGh3HDV7E2y/0ENewGpjp+i7w1pRwVL0JwpsGnDGU
dayqCC+5okoftf81ysmWFvFcV/PyI/7vZs+g2P4ZBrtmrewM3ZZbTTpR11DbtN/4
Opp6l6lbh5ysYT077whoPOw8N3xWH9Bv4ksGi3DMJU2x9DbRJhJevvdLYbHeE47i
b854+TU9xhSRKzxdMNwwzel7rmsJx+NEAWaWiPWALNblSsjMz946N00QYSnXowJh
a21Pa9GP0ODlXYS+Am9DTVe73P4r2Q93k5eWMfQZh5te/g5pnJwDTZuEtVcd0wSC
6aH/EC12MhkzG9mJbhXZXTxdhGy+Jo75nAu3tU8BMY/arqCsjrEOcbN/or66mnG9
ninudKDqdU/x3cOzjNAqd+doK57MrL3qv7zoUcRkNtml9V3dGPVaBPTb9/iaa4Js
amB7vnB6UZAyF9KlQ/bvpmlGEGf77OM62JUMmRH45+GpvSltvZLadutKk/uEiLoo
XTh9JrkMi48+w/ZrK8mqwFn9szSTfD20riV5+YTnF2h0KX5mRbYZ8BGbFSJA1r6+
hPN3qsHQVxMvM0Cb2DR/ySyOwLdE+VRAN/nshnmZ+94ql/xdw1cyrYbObk+0DNsd
TtbtUfPLjOxTYfbp5atJG1gPtScKT3vCH3vF1w5n5hFsjfECUhkMJat/QmHOuiFG
IoXlWmFHHyo2m1dkDKFbtk6yxmAfaAB4msCR2ByYdFvKww4s9Q1O0mvcEqmtUGz/
Cc9Kt6Ep99txa+1iYSd9u7kdjcLmelbWPZoDLqFNxkpt+a6TDjOTmfoQvezol3kB
W8jCRhZMUEIVFVrIwkQdpfo9NKZwjZCRIU6AtRW5srnqXodaUKZG85tx+snkzLDh
7e5a9hyASNmDhA7IrLMlgEsiF28zS6u9HcHzcM6joxYJGeBFcZUb5eG4h9JKJoqt
mPWPDMO9ACi0g5gvf1Lk4l7kCROqYFR7KXSM3wd9U3YNncGSuvbFU0NRGzukrSjk
Ymfw2r0qBBCRlBPszkT2ihfKHSRlHI56SAnrbtKAY+lVufuHWSdqs/8k1jrhmN7w
SKmp+wmsXmYXVqTLytiSTzrD0G1hpC7OGCL+28uhBm2Y1cHdNHpAKkpD5MQMP6gE
y4lSXF5XNk3gT7Jvr3YxUZbTCO2bsvoP0C7smB67WM4O/BNw/6c7A4xUEzg6ApdZ
6Bc7YGNEK3llwPfi2q/PfL8MQa1xHpe8cgWz0pFYCuJ/uA2rRPtmW7nY4H+TrE4O
u4p56BtIrtz6SEawrzBGpbz2M/Een7Rq7+ITpaOQIUybwTk2hOxqE6w/3egLuxvQ
A5ec75osR0wvLgyMZTTjdwsBsm/73DzAC8XJmAg19diaFHDzQGnGKd4QJuN/u0KR
5DG2u6GZ8kt7jhBIjWC3v6Ke61gwdyEUXHhltJ2LQyIRkKxz1hbCA/THunMG0S2Z
O+Duu8DhFthqezT42htYOZCKjxp9sPyn4Xy2fKqbTphstAZMLhtL0oQmY1G10AKY
jBdFzSy0pg0U6aPNaJZgzil/CRkU2EHvckZqkweNSejCht7CfHG1cz+tFax0Jv4+
mM8a2uYWpa46sofhODctUjRmGOsJR8e/dO/sOzqhT4nm7tTvEXLS3Qtq/J3kX3VL
44+bY452ntOZgmeCzi7ytKj7ldZQ5izWXo1y9+I5xI8Em/WsBxjrfO9KZI6TAo7j
DB891KAYKXE9tyFQ7wK6BXZHXel2DBSvIEhhPHUtlFQuSZs1DRc6Q+RDDHyUSAoe
WO2Gl2efY54KBPnw5vpToKp14R7Juye/r+f1Ejz8TCN6kEG154ad7mZUqJEIIXdu
abKfjuB1Jl9NMI5yNDMCbrKw0SkPH18y8eZ2d5yC+UnWKU9IyYU0yZViGKRIA9E0
+1qv1HskBt/pw0K4putvF0uuHWUgV9+cVr19xMJBWj0Nk1T+kHqY7krERgNYv286
4ADOmC90m+xuTssH8aZj3Kw3ztmErbBE4S9/zkWkR6l3zrk1Ivg16xoR4o/qJO2F
FtxmU4ZmBmbc5o8VZsr9Ndxo3z4smh04foeuZ708ZS2VtbNt6ZHHrcRPcQqF3eyQ
lReBUk2rl2IoB9y4DCDS9fGYcOVnaeDSB2DFUIbXVdkS8PKmiPgJZovFFyciTL+K
XqtqTVrsXg3jQYpvIRJQYly3Ook8IkcFhBOIU20t72z4yMrxiNf+gdwVZDsB0Kzy
UQdK6LWRk4KRGL8rtQKUtHeNpC/uM6YSfhjTHOxCWqb5LBipbRXCAoTaNDQhSdKb
474+Kv7oRYuDaBJV5nuQsngqAaG+Mz7kOcYB7lv4x2/bdKTjWS05uy3QgsJSdFkn
wmdIXFXA9uObN2HGWUCt6IiWfIIAgVXZuPLFX5BHmyqDi/IpDIfWF+Ida8L7F+E6
v2KJ7hhI7x8SjwYVG6aERjK4l/H5EtaflFxShy9NtS2Usp0d4o8sc9urcJ4qON64
xFG3ztvCU7HqvqVJZ2hSNe9xYCVsa1eqfdlM6hoUO5ys4BdyeiDWAy13nsasfbQZ
TCqs46bR7X3BX0F11FLImWDiYn96MKPv1J/rKBWrMjw0pv2hTNM4G2b2tduQ8fPV
URxv2yC9iTv/KCzj313A9p4CRS5ef4Vd7wtc4aEX1QdVNEQ7nZbkgIDz/faij6fA
DNatele86kXv6MFigfJPgQoSY4jLVXwLRo9D0CXp+tnq3sbbZ+CanbPLu5YS0ZI8
XYReLzGS4XZbwSoqwzW1+l1GDywKwHwgNLpsN/mbYmXybRRdWXMDy1YoADk7iLy4
4Tu7ZwXqHBrduKFBQvPbgqmdFzfW0WqLiV5ZcRK9QYx39en7UDHicCEE18A4AJ9L
pBevyh4SevmIloDQRPHbHNePKbBDXS3VsvNUK7tPefRKVbGfRJPRBCS+GHgGdeSk
3Eak7SoTsdWgZKcLqhZMV44Q5g/ebSGHZWyut2CbdwWlmlOpPuWmTW1pCNohIMYd
aEhgG2usvmCjqdqGizoqIgMgoBv3og35wnC9uqVjZiVlmyijq7ZbPdFOumz2jzjj
cEekTCWyI1Xn0/PA26YkCsN9odiSLZhWV5e+M4KC/e4pFdfuAEBEP+tFWDMRmmIz
wtiy1DtleM456ZdmrzGP/fwVUeExSC1keL3VZkh449R1714RnRrh8wzgoQlgFqfg
MR9ytozarZGh8ujzlgf7v9Y1t9QQeBoGsUIn7SriUo/Vn15oDGBSCmNZ1yacB2Sx
rpxwywQAUDhDENw6nqB44hwqZkjp5LcQgDnBIblrsczEyOUGY+B3LKKvR7PWFo/q
JjI9dPPKcs/EKqyq5GFLP6qz14kO4GpuG5IwWja0wJWu9YUqmb4cVad0JiTsnBaE
YZz//DzyuEoVrtJ2WFN4GISjYf2oWU6xPMRrahLRr99bUS5g2Qan/mKLjn+q7235
FrrRlkKAXIh/bCrafjQ7gPOcz/0QTHUcLcoU90sQ4khgqhspIU4boC7yKNFn/Y1A
CZ6QkWe0qlQVzDKN71+zo1yW8Ci5W901K/enkRxIhncAyUkqPYiKLGbZcm3nDYyd
3Br0r9C6JJjOgUCoDbA1LjlOIizFQrmX4lRzuCrWOcQXPY3Wh6dUknZsmncL4xKh
h+jH2G+E3ulIeHZ+396dHgnLVHPzwYze1NSpxnyQWlLZsF4PiLj96cFo0udFrQSO
/SbFtHjpG6fQ8iYM7pc2HyRh14QtxJvuvKXJDPe5gIQpbBWfoySNDuNPQSS2R8I3
wJ1p40qg3jIWl3jTrfOHAQbX28/isca69Vh9jUKYeK9RCJHkXXLvx2OHlgJGDMe6
59XdPrRH/XSYJk1mVBSTn9ZUhyfQmUjgxNk7/d8EpHOveo5jdlJJT4Cv8+nizbtk
H9vvuSLfyejb80MpRen8AnmezMpfRyOrJ6UHxsp6kUrsiXFYcLT32+PSEHLeoP91
iekx1SQya0ZyLg6KT7CCppMH1UPw8o41+oBNa1am1D87PduKO6KJlaHZZRSaha6f
m72ye1JrnLaXH51pIzi2LggQbXdQURwQ7NvpnGam1HlrIu9K5DupE4Do1h/sKr17
rDCsmVkRmx0ajOQ9HKmRWNqMiBEM/QM5nmCuD6wAASgpHJljhGcFD3iJhX0eayFo
eFvFI8lmgMmir/5AhX7aoQI2zhI+Pi5iyWmdXuR8nflBU2eusuCCGyHah5bqb06n
dKOnJYWPJr5079m69Sxe/vNFP4TT0AXbeY8EqZMTs13x77+L6uqy0ew8aTeeaU/B
mudLz+ohGaI8CDzs1z7VIpRMMU9g6D47ASp7aniKBS1/I3wScma75WAVGHFqafCf
TyCJhAAOPlRdUxeYGs01VUMhmuPLgOUK/MG3eS08XbAe51qhmUQU2L139o9pWlEx
hYzJHZJMisCJtWq9VHnowdVTZ56G/txdl3a/X4l7U4eaghcOB6x4YzAFMMTIpItE
LDU+h0iXWyY4nWMXEuGAx58iqEVohPgij76m2UDGHyYYyfa0JFI3WXvPZaUyRFGo
MVOg+Gly7trAcK+uSloIHKbxyg5+GvgcQMLVSJFWoFK/HYOtZ5FWCIB6jt2gNaT8
5mq0ibFUTtkfvm7/kmuvUSPdO4Qel6xHqCWYLfAC1b2yJUt4laKCpIHA+mi3vMnS
CVUGqEilw9HqBxONDmkkXlEGXsk+6Fk0Z64gU2+GgTeWkOJPMjN+P/dMqJxbbcPe
t86++W2jmrkfR4ZFJWrzW9m55dAa1t9YBIZ3QQXChUzr7anHg3lnIpabYq06oktl
FQmfVKkcdu7FZbPovJ7K7Ryb2fQupy+UIM457V22a5KZNML+M1i6AL3yRlIKB/Hm
Xnpxw31yArCQ286EGcgm2VK3iYX4C23IQIGrCvhULqsrwTZtxv6Glq0omXwRvrGo
s1YZsZ5b9O5jUhbcrUvvrm2XMGk3cE3G+MMcDn8IRcs0Jnecs+EXttyeNwZGP3+a
7BWVkPrCvX9LfOECfjx8r/FhJafEit+a7BR1XH2Z6Sdb3T2ZtxEg9aEbMRC4GRYm
Ycb+UpWH4/nA4A7IgELq6mmZk07hMBo64oB+nOLOZW+2EyhYJFe34QfK1xIsJ4By
vLlkJ5eTNlf61u5tkayXefvuuQ1gZhLgrzOio2oVWeiGDptEgFPix79bwuAszSO+
tUOk2XBOlKBcF9ExPSAkeF4hbBUcyNKWcSNZ5YbIB7zJifOmupe88jTYj4v2pCFL
qvB80AQE60G6nNKmblcuENlhKMYlFPaHuHMVyC/5IZWb064Ux/YvFwKRjqPL3bAu
R/mwabLAeDx/xlNQqgUHREmN6NNy/sRUEScIUT988Yb8vqd54jgn4oTnyzfL3S6j
hckz1Ht1YnKLxMSdtzo2hn9jbvxFmZXSyN9YYqL0B7l+dYcCsBnboJEnMxgm/biu
ToxBgyz3eKu6BFFhOmL0+z99nssovBYemZAeXN5yjVhT+zs9wz3bQl9DNZM5DbUO
vHnIYvY8et9gt0Hb8g0dKwMJT9JeeshN7gEsfKm6RhSFVwcudrYpkInJ7p4i7Cnx
IX2Z0hfOybXjR1wcdNNLRJejqNPFd5oKhskmjs2LIM/8WNJ36IZaGj2XT5kLmyHp
UGmYbTVOIbfasKjhzj78ZiwWFzFwYuV38rhLEUs5PQ81SxYoBB+zKXFMoFrtwkIP
oG3Xqa76414Jz09rvh++OV78dRQ9avsLIWlGinIp5DUVsHl1suFP4wG1dpSFwU3E
s+zi/1Lud+hcdyYP2UI7cDETgxEFlzJm4yWvPLVhLHxk70NgwWc/FBxu9sIW9SB1
lHJYfoRSQnMMli6V+Pv+D6setL/TwNAqJWL4dUgB4AZDcCmR/i96Tbn7Zf0XFZTm
xznkFvKvgXUmPsYmZsUdFdeoCQOjv6SvJ/ADwJNsRSrXX8ZeOAxeLav81Tg916mq
8bS4TpeRu4yXXc/ea8WF2Qmzl3E0XamrTcuGe9gk0MQnYiunFaPsU2ztIPNh4dZ/
Z9ztrp251KNMDb1OBD1L6tiExw8AjVAWs2p5Ln+ajjqwcRRW3tpm4GiyNT7aB50A
WsR5a59IjNCk033VDBdt22fGaf20D7BOrVKkGjZSM/3fIlYXhFQ3zwR4qX9Kp26E
rjbrU8Zen4ZFGQpGsXqQIySdKeUoYTcQ22wCw/mYBNQFUpSTRJVHfTX/p+zWF6VK
VOJ15tYtFvs9z0cjUzcR3/Eefo8xAFx/rRKhB6Pjurvfb8VXVVQoERaXOcGtPSvc
010H9EucMEgOUWzrUr+Cyn4xfV4LPeALNsMLRKQQzYP9xhpT15yY9dxcjLRpigqp
KTtTWLdUmszXDN9mk1c3a75Qt+dvT6YGNWmJl+pfm8imVa0jrf0lC6eeMjBhxUgI
lngU20uXdApU5QxOqlrBey3tPc+MTaKBns7vvSf6xnXXd7o9/SpGiH1alppbU2NX
V0TxPfCAzmZ5W8gmNLte91WWl1JAYDNoFDOFYuYNVnMKv5QzzGc6L2q6SGRkQQ0P
LJhaok6DfcVYZqvMIfkaTIqdUdx5BOcYz5MQnxbtrutLuGGmSAmOmpF2o5uZaqNQ
++FkZOMwOAQb6HPIIrJW9FyubQhJd8kXG/ePuExjJngdLJlz43MBTMrmh2PbzJbR
GgtO62UzSO4CG4Fb/7/Eq2gD8zr1E+LsBUnh67FtSnt00Rd5grLDBKcjfxxf+J22
AcYuKP4TK97KjuBFj22XfoC6DnTsdNHri44Bi4NMcCNm/aier+S2NKp26AEMfvWV
9vSh0hBrvpZufy62rfTZWqVRIo/TW48UwiZ2yKaexhpSFgSMXhn9eMu+A4JEyWQL
QlYlO9+7fPbmjlHn505YU77Wh5WxjdmZZWov4oVbXKmllCMmZdNRkbVqTMBWJG40
YDz08FzPvJp1zBZhRlQQltbJBQNUu7XC98dq1m/CeORs99+HhvvR2/qA4huASS/D
HtrAcd4xGmFmF3gWHh5w2TbLHBLFyBNTG4hPtuOco5WJ2RhhOMGnLxzjDYNuPcbn
vbaC+jxY0KHXjFIhYeXulA/uoGo+E/lV0GRvnrHN9GuLm7DPd6P2YaXmYFKQwED6
OjGmwSN3T8XNhayCbO4fxq9aRDx8+VZMtYJbD+Fh1IOGkc1hNpWIPUSYWsCMuXN/
qzkgxtgVCFdgTcUHq/sFiEpOXpNRixj3R51SQ1hrOjcLE9T7hKtEebEldbbHiUqI
5duGh4/6wfM7Hhxaf8WRuvGj+jGJtFsRd2h81E6J18Vxc+leQMrdRNb73oVCzEkF
9uNYUqtvJsF8e1VRl3AipalIhgDM0VDR446FzkONr5vHtu4BUoLMkkiXweONrD6+
BU3FDU/sc26/W/brABBTgluoSV+DrmpVj8qHST0ieTJyGMhnOhP/ZIjAKgKNW5DA
BOpXCPgLGFuii/EeL6vdkmfgOGaBJGdZy6kKhXqdQD/R/Iy+Le1UrgBU7DVBp86y
CgKak/Cdo21iy+As+M9FLddytuJi5EvDa/jwHihDC8klalZBD1Ii5DSYFEMYFBuQ
l6mdiDu4L89fwbbj/SIYjzMMSl5Txwfho+kvwuXHkpcNMEOWEOu2kPdmAM9C2fcN
VXNnhX2h9VqD0/YRK06lWx9/616hGSXPqrJKqbAY5xVI8M0bJZfvwc2tJ5HrOV2e
jmPJoLOX8rIkFCaMWSRHOUlLlnlnc5YlLsgtZQJ2iySrAB7J2uqMXZSgGjNWHz4u
4FyjeCCSUK49rpworAf4TGiEzemRUolynYiGcecD5hAXETMZMC0VNNwTkKNx4Ewt
+AvTNI+5hy6APGSU4qsco0hOKpXPiRi36yr1pgTuxqfvv7TNsyJ94hN3oep6CWaa
muop0xY/1zVanwCWgbeQEkedLY/YBFSplm7EB8Wyr5tK+O77badB+/YRYS8JbshL
PaAtZxIM7IAyGRyhYduZSEhqut4mm7+YkJ40b2W+BEnsxFE+5FpLzLDVx041Yknf
OpYxB+ZgnMNfP3QzgUyLDY33nInP6tjmcF+lBfgdVndXEXEl9tT24NKqrVgaxGuC
K226DbW/ux4w6iK7eBtS8MLBi+n6WCm3FQVX58b64cqkdKwo2ok7c0reTwziqQY+
GaRAZv9VAKBACJmotUlbVLjEIS7ckJFSvOxTmfJsH8tmdNa0W/qpA0XiVpMhcDXK
8dcVm2RXH05Do2j9RwCkKGf3wh9tFSgZzGwH8bRZL+3p8dM/gHhN9c0en3nFcNAZ
i0vEVq1y+WFlPndEjC3tcJFnMDh95G8JkoQG2Bh26AB/1P7mvWls0vgEud4yeCTu
feW7X87MddXsy7CFwl69i4MK6mT+//+ocljX8TJaCKDw+35zUOoJiGuIuF6yGTAH
Cyb36cf2hg4DgG8PT21gKj9fAyppuPUbGoYoYMm7vYGLoeVsXRisoHWdTDO4GMZa
VnuAie6RAZRRR/3VsgqiDxDmBEAd1JxFDMhD/xJ5ez70XO0FKYpJVei+dDERTPGP
iaKMq1mjYSaah2ZR8ddnlFDB2RwYkmujdsYIOro0x7ippxNX5+bPYMB8aHIf5lca
n6GK5tugxLQo9bulEGnb/wE8+irr71One2sN+UO2OM5gsyIZgbUdRIN/hFDAMh25
hO60EEJPyrllnQbO8iQWHkNXiH6I5tO30OSKsqYqe3fGPFvUr04HgF94cA7LUnG9
vY2LSNSoRk29ziQNZpzY0IHJVaxJBs+gvD9FauqQ7IsBxDC230H0YJ1WhvA1AXXX
ax44a+L+Dyr+Q9oQ3HhqYgCmrpL1uLOM2qS6R06qUdkPDdx8phdhvSBWj2XKF04N
fmTCEFW/SThP+fBNpNmHQmJM2fsvEjrf7hIo/U1GfYp0DMMgPj/BzLJCm4cAlhDz
4FkF6yhKZSCgt81mnlkjxW6SgaLH51xnLCVTt07SdEFcrIdqMKUfxLIixHesEWyv
jblM1Y7YwR5TmjTBcgOFpKJkNyvyuMoPXyPQIZcB4H0qRUSuLluFPSKO8xNS+5S2
Lkehgvh8lUa6AdFy5DCACbpkvVp1xeyzxD3KvxNu4FFeZjC+PgkwEp49u2hk2Njy
a06VMdK1ozO5uLPvh/+asI7SLWEr0p0VF510/VkvXMcbZiX+nP/NsYp/gGPvd2kG
y258DddE9oNBh3PwlMibzQJgZi5ZfIiMU35Ff0hbVKRPOYttfogGi9SYQ9ok9FTz
cXJdwzrbSksxNs9Ws7ckUHz6Xt3RHBfQxVNZUKaqi5vWkbULmnacHyhcRZiIxBqs
jXjDZwjwF+Dr2iG4Gb8qzpGDbupy/xnbMz2e8iPvaFQROpnf1VwCrNL3KpxF2tIZ
k7KtPOICxrdL2uIX2HqqQ3JM/e63C2QoaiKdyFGO0D2XvWypCbcZ0U+A9gAaZK3P
fBfM0iT6hbmaLR3vV+UkHBg4ZMbvaIjw+od41SC5FQ0JjGBwzrFiTr1FerBJXOHH
cVtRKZ0TxTLEDJgPbMiP5BW9qqhIRDVpoLc/vp3Q4hb2VtbBIujE4x+VmbjU+sC8
O0HOtBLn4Da1sFB8CMcS4uPd193jwIkYg14jVWWAEP2xN+YVbB9PlKcWNijESEXr
qVBVVREKHXU4nEhF5tf4ump/0mYapao59fFCij9jbYTPRb52evgoK3Sdlt8XGVG2
JIHxYaqN/e9z1gn7OWA1rg/3+0WC4JHk2UT4isuEoLNA/kcWf73j8hCM8E//BZwl
D8uE3a30vc/rkD9OvK1HpQKQEUEMLGx247W7x5iiCFdKY7tbOKJUm7z0P8E+k+6K
uPt2jzjc4bfse0QzvMZl+5Xn4F99Z9RyRTJPFhol7K0LwREEDOIAyg1MqeEtrvr2
z9CYmIehaJRfSnh7RuCxFlqv7GkVm9/CHAMhOE8nSYveKG9T8J29vAy41YxJRAez
PNNs54owZW61WjsUpbIUSdHCE5MdADjhTu9gr9RHuaT9mNHNcWuR8SR1RSPhMUn3
yzVnIFDVTQiP0qqe2LKZOji8qtQ5VDyFHLOqbRdgV9NeDBmYYuWffS0hlxuCYkRn
DqVRf89/y2m4Q1FiiYhyP0DS0XwUo42xGM6IMlabSvxw9MC3DUKPXVCTHiv6cUjU
uYSZkSHpE06C8YA/HJL46Ljj5ApwqCm6cEHGRe3ee8Q1tvgdF8+D9cPwx5pmDPM8
K1QNkdceWm2kf87UI+EtlEjDwmeMdlp47HfIMskqrqvBQ3SGkjMWXv8WRo8Fghmp
TjJbBU2PJrjWRp7Ouf0QH1AlTB2BWXrGcxf8MWbeO0oGe8naST1kjBMbiHuAnZii
71kSC3U/0ZokwF5hUbKRVVk5RWcF3DsnhdaM5+KS7yHTUqBsOrm11uONeE9X1OnY
VRDmgza4wXLxbzf30qZWuR2WRaw0zH3ijKj5I2N84iSRjckhLP1CuV5pdXlwrAuA
lD2XyLPfzHnvvNox879XTkBheYB6GQpdmEcFrERXuTlM++y6X/ChoIib/iXbcRZ8
T/q77hUsORLM3uRJnw/kl8Dkbx2ntw1+UESQDNU820OSQYsjpwMofDAgu1zCgehe
/kbAAB18ng965KpbgZT0cZ81zb7BwaP8gf003lcTjaOj11brP6IdPNQKCZQGyaNr
dKGOLrtNdhiNv/RnBs6sAEjt+ROd4BEEtuipCLz1kumQztewOrf+bU+qiNyhfgHr
a0vBNcS0AVRpfNyGJ++DJ8+NIrgpc/hsgGOEWfplbEmwpguylKjzZSYferW24E6S
7V4lGGc+ZIMutx/VpmGrbdl4MG6gjicfFNvtXl6disnB3hcUySJMGIVzYjIf0n8R
X9NghiQNj5fwRlZWyYrqm2fdqN1ZL9AY4qN1EHNxonfd/Jd2Zc7jFbrTy3f8YOld
JYJEFHodVAIJvGJawff64GtaZdktDpOex5JlJINuNdkvrul3Hj7wT059uTWgS4wm
SAiFCi5ziVsPBMywPbP1OFJxQ7jo4a/ONuoVJFvuhO37CMb5LaSuiCzLAz5OuVEV
RX3YrEkZ3Yopu6AwBvZGbNfMDP0QxLssvN0gu3r/ds8XtW8kXQsl+RCSPW5SC+ve
qiYJQgGdUAlTneeNdXFxVkgHz8fBurnY3czdjqb1gXGtUD+1m2lA8EAtVeX/LzeW
AFROlunHJ+hdRuYsQLDsOq+5knGdEIfeeZlbGS7VInbmB15orXOOTDroA52Shc/m
ZIqBhR3w0z02BDWyQJgoKBL3WOsvH7kzo1oAjMQJlz8A4KM6/NJvTFMnpJclwUu6
1iXN/tgZcsrsFZe6z0HlPcgw2yQ2cEyyAHkJxpMdjUWNqsbZIHEQv60tz7NNTNO/
t30cle2pRxRtWspdqPhdWOuqiYxxCU8JfW/aZ+oZDDCaFtHxuH15sYrDqMhYFHPC
jR/DX7BCGjhWZWO4bkEfMVU1DVbfSRjJF38nxjjKlOqEHHBcBZDxp4cHU3Wm/ipv
Z+8StLniA3a6HuENEedrG3YbJjfMxj+0nmqqgtkrQWOy++oagHJg9rKdEbe1QqYx
uox1Bx/zmvSOk3v6AbqjVttU0etdIXjiqPFHs4z0QCJJfIfnSF8eNboGOo/15jTW
8ZV5HpDekL3MZHr+pjwzoembdt0XQvD2zq2RFA0RBhI2RxdUm5wxTxOx8/ipVlPX
Dec0zOYtVkBhH9rty/noxdYVIJLETtobA9TCvQ7rO6nmSF2xYWZ9t9d/FKeuA8uG
vHYqFbPKr3GN3Hvx5IuZ7R0TcTUNEbRqa4FMGwlEWSUYmv7ZurEsNsdIcJ1ja0qq
gAePUgmEulPwzbpiuZpzwFL4LuDn21Y1p3qHi1yGq4fFfvJFE78ssP42YS0b7rEx
JBWNEG1xV/aiW9b41Hvya1pxyWW/bg5MsskNWWKoGfY7++yJH4mjUThEqm5+WkNr
G3dagE+F/vq1y6/Ikh7TnghKdrGao3JX9HbuywuThLGClFCkUx3vKid2PMjLNuu6
0wUo6BIaCDkUh3BEMvZ9Xrnggm7xUVpXBtD9lcSv5WmQtFTvFF2j64KX1qniW8m6
4WXYe72IfYdwt8Uiouc4QITbKKFEn8ir4cA5O0sBdu+GBVH9FDXgHZdvj6Q6AG5q
D9G/c8WkCCo7GNvABb9usRB2sfjzPzu4oK0CTl+j6Kcb6soIS4lcSySVfxWoQi0o
JSAKKhRH0WJ6RDHuNPRdCSze99u0Ln4Jijepu/S/4bQnvTTzllU34n7FJQQDakm3
Ou3DCSWeGeU6NVnOiW9pXW43n19Y6cbsRT0kszkB7g5iuO9E/6DGuYrBzZleUIv6
DrDoaGckUQa7fVVd6REDx4MDmzDU2Iv4JwqQzW0wstc7fyxIRg/jaOewr7yV6Ax6
H3lnTmL+3kvz4Xjd1ju/egehzkR55CJkcy6NxXrc8bo/AtDZQe7zSQV29PQZW2sR
koRAEsF0XgWd9RFIjR5yU59p+0CvHaiPxX0D/NOLgGE1K5lGM7gzsnU7fxwX5Kxw
hCoR5Hl6IV6LphC6jLQpF7KZPx3PbBd6epXySugC47o3S6Fb9ax3d/hAJRmKIYB1
XtLIdegVrWNLwG6M11MMyZp/uayNb2WxV9itaFBnsD/VtnL5A+X94YgXyPfSF0kH
fBEeO4xtDWVZLJptMNSi4voHjT4suQXxfEXol4CXetbfuyOcAJ5mcCiLfUNz89JZ
4pu833x3R4nGFS9E/N3P4Hkq5FB/sv9lCozPj7rlNXItyQ9ePLlIKtdI6LenGml8
qDFbZuyUieFXGcQV84kOD86jIXuXHv3yKysE1PXVs+crCDN3TGofM952hWdOAe4X
bLF4YtfeTOIeOk5zlMVbAHQs8xUr3dDreCNPTF/tffC4d9+HzDx68PN1gWGOmIXx
W3oWruAeRoBEKqYnJ8Ns6DrTd1l6eaYDS0rhk51alsV8eyb1ClKAYmwqGzdI1zr4
i20A5C5jnXuyZ2zMJJJPX9nmWwze5C6zgg5Znfs0gr9floQXyMk7dtDr2LEcrhBu
dIqF+amiNJJ+BrYvFB+osjWLtZM8iZYP33uIq6bGZVl968z21c56lN04ecAIJSce
FtvfLn/JHUoaRFN0QWx8tNAPsP3eUCTvM4atPClUaJg0p5mgfnsHc56JDSM58RNz
ZWH774sbP6sIjt3XTD2rOFCKQd7mlyGOIgdD7JWqyd9o5vQ/5yEZ8LjW9EkRKFzM
J1vJlHgaMFeCfgPGH2X7QtWRqQRdOTwCf2X7rT8bu7k+QwvZGkrmHT0tGNzZIuWm
thY3aUXX9LriMBdYZ0AFa+2A8tASKM0FLr0oq5GuLAlElvOxlcIKF+VrMzqcXHo5
BokJZL0l7LrafWcWr6L7EpLvhh4GAd7BWvFfkBv8ko2HYgIyrN17Kc8C5BtRTJea
A/oHBucchzbN9g8f7EF7vKvVqpTI0/haYy43omPV+bSN1DlgQ+EFPuhi2ooXVY1K
HxK+lyN9OdAwcg5wun9Zk7WONmziYWYxNbiZd19lEF2y5EtwLCA6ZCo0RzEkpztI
T3Y1E1t1GuQf2qZyB1/QEcZKYz6MP2+JSfItQ2oOHpgRGxtpH/zdtzdPNhCJNZfg
eOVSPZxG3QnN2+m5TmFbNuPJE+egHwDpzDy4KcAPu/JnJFaysH4atlxytGv3EstG
3iS+cVUXyfgKhy45slFGczxYKPc0rAHqi2uA4IHRZdS+zlfu3AZCwRMWwLSu84Vm
eQx1EpIYWW0aLr+SQ5RrKiqmfYyfXKv8cPf8GZV+S6NIcZOcXNHrCVr3hmILaQCg
YpPGzIdwVQ1wqh9scqZdolR28N5p3qCLYUqI5kyRIXbqMGjJEdZFW3pLMeaNpC37
RC1qXJ/dFTtSUw3QjxzW/id03CWj3gAcRIFXbYwDK5hT2IvYgyFDGMYQ7LRsjlsm
EN+uaLqfYVgdlDRdtCYqIy8yIdtLZt2AGtSIRp513pfrzQvtKg30CeMJIISau58R
LreqF1BqvujCSnOU2+nteYv5otZxDUmuZ8SPs/EP5naSGDFgM/3j1oExY1pRdnN3
KX/39VFFjSnP90R+8Y5bGhE/a96W8NWGZ+xhYetLq01wCPmUfQWpK/DKITxUzKXK
gb3M+/NaSrYhCHIiBFQIioOTKYj/HH9ri7OLLSkWiXyg1D/QT8QSoWsXC7EGmI8d
ANYtlPN5j0dIls3+XwNeuW9jMnC/Ru0nQRAXOdVPa27fqc9gDDhk7M0ZjyeOzIeu
R9A3Hb/oMWMMmVzak9a3p+tvzsFn6qATZLvGPFY+mohDI59gvu0Ser4q9PMJcJ4W
eUooNS9FqTwKBjSgQ7Gl57+G2qLIFqaxiQjIm+2IQbYFInfLlHDJk+l9Jz9rXzBE
pdPxFJeUEyAIZeLJLwaXHMTIayhfDQZxm+wYT1Yu8rnHrdD1/RO6XfOQ1jrpuKRO
71oIQnapLb93Mac6Mlwx8dh8h7hmQrZfei9NzDegEn4MCZMn/wYp+jHQmY+jQzyb
DJyISBaNqmHhfeFmOtxhbBCENqHI3tnwC1SorbxHT+q2dCyyTBct4RzWKGnXAHNH
znWSztE38dHe/+7McKabsQmXSLTwkHvtkVgqlyq5ENOyMXhdJvmLNUFmiSng4i6J
QOtUKwVt11Itf0v9ts94vkUiGRixlxQ7gLc+x/7aRqa9BJAexxfHgQureHJuZN79
1ViCl5WHgPIfekTAoTI+xVGk2lOZ35Dza2kJ2o7g6wzamBv0J32cSUzTkV8nUR3B
eReq8le35HVH89epSi9Ocjlagi3l6vqljPcU/g9ncd+NJAOOwV7yXAgdAjmo8Tg1
2C9W0SvhrFr5zKZYDVPXefmvrsmHYO4BkneTwH0cQwvaw0+sJwHQucBJyc/o62b1
tbqL9x9u3QAdNNYDu4MclUZrSOXQ1SnkfQD4yfy4Csu0GpHN7rgZhMyYHQwtlAbw
IsiVRxjJvtxPZNAqrT+a2ry8sHYUbQVU+eWSUDRYNY72WYVipasI56bbfQVCfyEP
ld+yjCgKy5a2NzZspS/RRtm1e/Ndnoa4zL6kJd7BIQHp9u1Gmwx2Ayb8Zej/3sWb
KzhPqDih5NMxVOL+hbhAqR25OAmV2r9AdbMHAi3ELJiqtbJinVkpZMer9JGEf/XG
6BwB3mUVFDoDC2as2F7TrFMiXKmvU8uaD9jmTI9TH23WDhmBZ/NJz476hnX1gb8F
9TIduAFBEtQsBY7EE5IHpFojOMiiYTsCDgfZ81bqjnHOg/1Bgb4/jdUGrjGE44KS
nmvuqwlhzC1/FSb3m+JDzPb+92os9Y1xJKjmNw0tz4HwYRtADJOl+WN0OahZSjrL
kEqIzB8oVptqVuyqg3j6KI0T6QmbUa6YzXld5/9MGyS9v8j+3rWufISFV9qSzxlM
N5on0BKk0HTAHaHb/RMpitV3tg7W3Ad7HvGY9Rf2PTFxuYkvmkb1z48Viinbav6g
cGICWFesIdx/tm8mYaX8bpcMv57l2kYGiMuFshuIbjBgT5bcxToHB1Of38+Cnxqh
MAeOfy2g56RdI7DAjzbuiLXbH+37spwVsft/0IvXwQhYh+yFpbMfzJQUjYMXcbXn
AyMfs/ysc++1GyjMAzPvUlrb3WwsvUTJxY3mh8nfhnhIpljq5HeFpKlvvYcMuCMD
d+W7cjGNnnDkwaMZSqtGVnev9CfDAnpGtFqffkMjVZ9kNTVLCXE3GIbaYhKhrV+q
JN2qVMDnZQROfrx041vpLYcYcxjyHeD2sGS2pGy5g5/qJayfeR9ewIvnJiFGrJJJ
a/CCqe2/J7bwC+VObwRcf8n9YxPNFwnobSAZ7oT2T3CrZqHKb+hD176KqKouYzEU
hdHjHmj1O40l26VdlaYuRT6N81yp+AZqMVZNFdRB3veufQk8Zgp4/PjUCG6Sqr3O
ESch7Ca71BOoGwvQC8t7uG1THgcbWI9dm5T0tofDGlYJqCY62L1FVWxKnyq3TKUg
EDaSnclmKRmaIdlXyuzWPPvmqmuUDnXwRSSG0TDCGGtRef75JQwCuUd5ywrwrVbW
uWDtEo4hKaPmsGe7W8YNP9n/6NazEHVpOtvL4GkQYDh2CByObXrNc376SFDkHbXD
3NqvRqka0yh8TJosuymGGWtvFuSd58hSRlvZOoHRf2b0h0QJNyDwbmiX46mCH+2L
OjS1gZ2B+zEewElHFqy4Uamk8XkQOQxwPOR7940i7ZllpRsxyVAqi2npNBoQaTXK
9/h0kh5ZYXP6kurzW4a1HhIxOXFkG4oGw5t7kK0S5fRIzRYXgKcV6aQwlYtt9Im+
Xx34M5yOfBH7CedPqt1BYvtX0fF85SDZ4vjDK1+NCR1ExZN6rYpbkO/si50HHvqV
WLUGZvzn+ZOoF4kKkYNolrils6rn0b30MjmrZQaMYpsSwTiRozdbOXD94ZEU8oRU
m2Gw+vsOxVPVhq33hTZSLs4OCts7InJHm6oLuI3IbxVsG2lR/VtENWGutOqQ1A/I
BZpMCKfphVAYiVLllUzmlOCkxx1QoIMIWqhEHuO7NMr4qzWR4WHQeJpE4Tym5DfU
q9+o0sp25NqjknDmQ1wPCsculLaSXPNtDzrRd88tQb5PHNyuIGvXvo1NMX1eLp95
cDxLI1lpLB42PHntDHiOXF5labzQfey4aBnhJOX2YBxTyy8Nf7tuf5OrDZ5NPmxN
Q+sDmVcMI3j6VIBuoJKcxslPQmDUSYcypMW8qc8AMdC96NYgcyEIfGIvFg9JNf6X
/HkSXu5DMpX4GHD//lANq/mDNY1PN0XKoOjXbcMzyAMFbvnIqbGrFt1IsqqXcF7Q
EXhMciv9R7WSa5GTSeGN4ixXdY5gKI1g5RY+zESRY2EM8xG+/f4xwWeXYrloB6hn
Az7MLyRgIKclAEx9TNNRzAQUxRxTJ9oW171f5JlmD8Fhe+3Q7RE7AgxgbZCJcBQf
nK6lIKC2uOE+dAx2TVI9cdYsCiwaQ7TZBjrF1WKl46sQxObrOcdYB2o/psDLdrpH
/6wg72CqEHtTD56HPbaviN80q68H5AXjSZ6etjFusoLrCBD5bWwSqZSQjR7D2agi
PHstTF5GyD9BiyUax7NyLxvqmM0THw/GyfaKdJ7U4mBXxGgdgdzJfMx/mKLDGMcJ
FSNixS0Ozf2jzHxjwpoEhA8/jXRsYH7DxnZ81RYq5ZCL3hwWLxVXmuscYmhoVWkF
+J+MFIQQTx95Ll8KuAoFVOsXsh9MPlW9Xee7MREkt+BzhdbL2mOOwonMqD3fTCK/
sWPU8zbNj+IC5442rPosyKTjOLy+RUjJ8Ss+/U+NUnGPCJkDYdBd8b8SNiKw/o4v
3Pe53dDaeC4GBcHwQUoJObEaB5zGuOO+/BXgg9HeTxmuriT4nT71XfsW5jBGBP3v
+FblzIT4g2enW3VEUEm+L41UgFlfN0q9vJLeqLjdtq2ukOEo4tep7hva1NyDPmxV
47GWvcKhwDfK+Q8h7kC+SO9329ssVYU1jtfmG8S0HDpPZ5D6xj9egtWHuU17zjym
iV62AmSAjxRhdZ+aJYdu3oErD18LWI2VdhgknEwT4O9SxCm1uEDGH4iFH4Jj/hPW
3H5U1HrW7zeQmA9T8s5kUXOztNJuEAJ20meZquFGRjMv6U0jXrzHdDOZDerQmVFr
VCkFeARviBb+RAcycnQt8o2jwGwE34wpDAkWmAr9PSh2MS+VE+QCD8blYXgUh4cL
ZlrlCLhmOcLZJHT7rBvl1tXJ4THUX8pcmyeDLDPJcHoD5WhXC+4APFjjKqsO/ZiM
2hutTMqp8g6RKpdJKc1x/NDnoF/e9Z/cxwp+g/riN3ALCpld3BcRQ7YQg8Vxo8mN
SzQkFohoR7JeqTAL0WSO4GHQn5oWOXw04EvaJj9YtZhC0uDm5kSrEuVw1IAMU2Kb
trMjEwod3HTChMqk46WhQQVDOEtlO7xq9ljmjxHT73An1v5g1NthQsg1KCFhMHc4
VoLKrAPt7m7/nNZ2fxCdGG3wN8YvbNbL9ufERXQhVTx9UjyChJ60OYGT+m5bUwOG
uT80n2Cvp34Zs+enUaQ572Q/URJP9eOIVZKsmlweonj7WONEYcJXiYucBgU4Hew1
hdXHD7nHwJiDyQ5nnUIG4k9R0AulsuJZM9RVLI/vi48zi5TZS2QH0WKewo9UhxuC
VWr8y0a5oflqF/KF+8P7iPy16xtw7CmQUxEjKJ/B5pExaQjAu5LYSODIxjt0Llbp
DZK6H7SGczetpt6kiCr7nd90BSudBLXYW0KUgAfV+NQyifGBWGX++G7W3O/agSlP
ILnzBaclHoeKeadJ+prKumEQYmOgMS86bb6DXLrgF8G+zQV9bxpqCoXzBMKptBsf
JHRhVsTFeGk2f5XlMb/ratJ81n7BDIKpfOiUjNoks9+ulepW69yNhCv3UrZAvKOJ
g2lYJfM1/3L+jM12EPD3HjfHzvDQ/5WFVDeeCnzehGlJRsNb4QsSvPTuhdCTrOPd
YleSgtah/dMt6CTq3OdkgtdKjwPTLEYJYTZeCzR3lnEBCCMJcHKYI/G7ZVIG5Tnq
2a5DB6Hyxcc45iJGwwkS9jauLL7Ks1I+isEASHDJekSKgH0bYr55T5yaQ0vGWqIT
/FZpPy/+vnPIBx6eZ2Oyf5U+cmgHN5KlJTDmn0VFgebQmO2/IraGwIz9kdgFCJJu
Yg35LYJTeT0etAvaXHlKz6iu50k+2YXzCYYrxfeWhiZ7HEIzDTJCMfAAIsMctCAQ
lCRrwKM5Fsj4Hb346htinqTO4cfSU/d9PvIEpW7QjAptzn3WSbBxsEHKzsvkXeX3
ziKR82j+EixjXurCBC+3VT2lEceHqUIzKxPDmplBzB1vnjT0dMRpzpcupI+fUcwN
eCvmOuTwbEhwM5wrafxQddkQVPwvK4+EoWFTr7hKjCjlYz87XGX8YPV6Y/LQqrm1
COyEvdJ1ImpFXGNi4+eL8aS23ok9z4KrrwdL30PdvEGYV1eM/WbjCyytXrm7+uxa
GVdLywMIWHG/UAQRc9GWmNikaaALq82YNKVJVr0nkBWp/HLNmWggaA3AtJCMY/Rk
717grVDETo5aLiS2GP2rTmTuRPGDdjphkFPxa5oj8nSbJ6BHY681o0MzW6ocBtgZ
tz5hBgtgWHUEUXQcJaR7vYuq8npUf7HhVTiTICXKNuJfChVEIXVk3vtjTcRYD2eM
aK0X60LVPVAetE0GToHT/Gq6ZKPQh310mTvUfRyWuY+GTh/FOZa+yB0d0Afq6S7h
P589sAYAgt+frZM00JK4VMBBylLfaM5gAtn1uh+kEE8alJbgPmIpA5xBtl2x0pKm
+dTgRn69JqPfiGL4PraZPwHtKWN8MdtWpyNGCgIdvpQsUK9HufmxL0FMnoSsAn5t
GAL2Vw/zI1qST6oi40SGV9IQYWn7tFPcnP7tPyr+xl2ut/lH1xD1L1h1aoFBRF6k
tY+htXUJh6/q1/PRYZb7VXwuW30+9nmpcB8Et2DqJQN0muDHQ0z7lp2W9r3LwWee
m6uCD2tYCuz1e5sE1Np7dNHC5mrjp1izijjsHcqwfU6ikw+SRt1IN07k5wmMzNfX
/6IltR+w9RLl9auwxAkIaBW6fd9ACuxJ0ab7qQGIBDv4h27AEzg7W5BWc0cRxpen
97UrMbTewXXZ7c4IiJHVZQOjIugVIlO748BUrnc12kFcND9zlyuzfy/Tc4D+vc9Z
6rcND71saoSK+O8NK6IswO+2PVJjvIJlq4DAvNftFEDsYPpUB3gDeRjqXyDaI9x7
JsnCLlq5uEk3CurRhzQsicXVB6eXMgmQm07SykTEu1fm1uO3hC7jNJPAw9dW2zXJ
iFSf1UHgVl+yRn7ogH4SBVaDIc3wYlSW5CSGkhboLhMczeOX+f2rCVvDPMbDQH/Q
RwRj1+Ro+OHQXxW00Xq/BmIGeznkWiqxuO1tO+tcLeFvWci1/Rm5FzaFEx6QbQo1
LZ9rbLu98JtGoOMRQUhx4LHF4mnUroK/ek74K+9G89DDDThWBFRtsCUu/9dRhBC1
j5pPWoLn8oEiCdbSGJOyW1RWViqhQTyqavAMPoMqWxDaMM5AYJZ/hYZbIguC/lXF
UZ7BSaW50naLU1jynN97ibIB27jAp+3U8Drdl1QtCVWzku3ZlKydiOUzI0VMA/bB
xWXpUsd5t/RzA3J8pSNclDm/5FI7Etw9NHmHg9jFhbPpigLdDNIXsJ0FmISnJxGN
srcLpeU/5d02vVBfvypyngOLWfkNbbxc7/Ex09NwQ9enPnRfmRDwKcu8VWnUVgmG
PxsdZFYfZHkK1kJskmUjxbj02q1N8MnfUSDSNH4KCxFFfRHJ5XQtQq2HO16WqO1U
SA5M8NoEkItUewljog5TzNRWeOKR2LJQ3tVGP5S26FUnB0NxCz3a2zBHZtfhDL3x
aZGDUgj8WTxhkeE4+95rdhECnQLUEtYpAHkU1SQEsX4OdF8MLBObCx/HmAT5jL0G
iCkcdt2oPMQC18Lj9Jhtxv8WEuU+4B4yYt4h/A5H4qIx3g1zdVtsAyrw5B0J/I2l
XXaXCGG2JMu6Ds7dB81vKf30ndD8KNCg4DFIl+tJtTpJE7Ot73eqr2L8Mpa/PeyP
rWiaPAEWfxSAC+SUi7tk2Q0JM6cbziGVc7hVoBZlRcNL3F8iW2bmJSSDqGMXq4ID
PL+fGfkhVPXSszSpyzxd+KgaoQOYRmtvyI4bOwolXfgMqotBKpxZ8xfCTFcohpS+
LssSIS8SAANDkp1MuqzCfNTZt/ZCaGZ3FFD50iNu1gYMobKt4/go0RJ/mXr+8Y0/
y2RTfWsNNl1J7l6AgEvRGTK8ccF11LIWacWwBXaLq8hR3wkJG+tyFv9wVP6KDv4D
2cfkiIO7QVNhWbvWZCGIK2unuWA8xCl0KIX5T8uBo6YaSh4LtGJdaMesyBnujdAb
+mW6rDnOhJnzzl61/MShVau5NQ8NthTIAu1/xmkAIWKjxS5+jrP4RlCIMTk3jd2R
LSZoou4f/7SA6dBTtmZG2d4UxJPbv9HWhP65kXLLoLqaOdyA23EgzIiwshbGHLi7
uUO4E1JDUO6TVE9w1F280BQskZ598iiDXpdEuLRNRsAhmYwljjVNDbHlz2nbh+60
cvGrL9R64sVoNZkS/Ry2198LfPDlX/2Lt4t4SgYSoZLJdVpiloFev88hVDt1xjUj
iqOk8TeM/ZEXh57alwiTHG/E26nZhMNmdiNJwFe2XwPdPZUWGbIA3DM2XUHRR5XG
REmXuQSP/ovIxWpOBRTXhqhzXzK8m8l9J5RIhTf9bcjQBu0AqkyHEFEUUZGGoV5L
Fmkx5nT2O3oJFpw803XWAJMB2lq2afPjMvS02dOmY0DSq0noqUzqI5bfP0+z+Dzf
it1PVZ3RZMMjxiWt9dPPe1OFRPb7px7TUKxaakUuvTrJYFLnvaCm3tPUabmaNgOy
AuwNSsY3e1TN4Fto5+1ArTk7PfKFs8VMzTKO7pNEESvZeGxaoUO/PhiTLxbHyxpL
k9/fu7e2OPP5j63nhVlC3Iop7V5P+gtbTW4+2nDNJfJRnB5Unt3nOLHYqmY0hUzG
K0zyP7z478K898wmAUSQevnTYPppbHNpBMJu44l9FAyKFbf0exUzLjdu8jwGUtma
C7aH5GVbq7BQbuiWcxI45l3Pd14zPxcQmGJMsswAUaiQSIUYCXnZ/aiE3IDJgPWa
iPzff/1nLclVrFc6AqXhIMQuDj/Ink0qG+QOv7SmMmySIahiTjQyL/Bacw9vdWch
vgOgckLDE/F88Ve5sHBTskt83xEYWePNP3uZD6jXhf0gemEp5qBTr3qrra9+1XbV
c5Ggd+IKZ6ction6dgAQ18Er0+5yzdkO7Om0U1lEWsA6qT5a6G63DXXCk/8Lf4Vj
DlclLpsfpTy9VaayCpShYv8PJNb77JTgLce400WgCRXteP8rfqRDL9r+RjIjCmdH
xGiiucfDZ/8NmPcyz871y+t07cl0hYO1WF3j4QKi8rwHf4fYuoq2qIUF9PL8hNlX
9eBI0K36/7mY1XTx+mcDeHzWaKbsNSKPNUX3LE30pCoyQr+KCo4VxEoX2+4mNc0R
JFjrWnKt5o/6/M4ejBU8kx2AELEYVH+g/HUYfuSfPfbGdeZ/RP9MBsmJ81poZosQ
+Wa6DrqkVvoZto3Sztx31yMqxPaJFTCRYT1F5rj7PfLnYF6z+idBTS8Sqyg60wwk
NdgNB8zVt66J5Fd5nU+0G56RwXHIBuH1ioePbIOCFsLu5NvaMC1eP9o5Ub0jo7aj
mT8QHfrqXdT754Eu9ndzseDHum6JiR8lPmUmOmvS8e/bvzvTHmm2+YuCkRUZTRht
HAaa1fqut8DEpXyO1PQ36yPIvbEJvtyt+Jclwyn+ajdcX6PLF0+UYh3aaLuKh29w
FfNteJs/t2Ukx1k6uI9OKzlPIwUwdC3d0vuBV4kumnWK87lt3s2oejIvId8tN59V
Ly9Qwkm6q5N1Bd7EOWXlyBH7SeHGfjrPsE5fr0w+ghoXxfYcGT23vXVGSYCSz5fN
EBphVK5/jhoc9FWSva8ASBtrOTrxY70sfm605ERv12PGdxf8jaBktXAJbmF7q7tQ
DB3IxR6lNh5Nm3maF+tHaKeq5+qp9eXFnydn+VRwoqvNF0zPoDjckeXqQB4oHURp
TXE+bInZzA19XD5hvLoQ1GO4OjJ1Eqfhz98e17pSM0/RmiqwJTTqSaXRCgGZJfhH
3g4VYObHtmz5dASPIrfg2ka+vcoIgnTwYgqU1mhLJucLpExBr1gUbeXAa7N9sA2K
77NMEQxkz+CAi78DIEKbMeE7aiKwAm7U+Gi063rTIGGSvtt7z/oPjdoAE5NeLTxj
XyzOqpALrHvmCaAAyxJ0V4aMO7SFsxG77TPKGvba93K5BbSJYysGu11UM/doKYm0
c7lFuIZ9ICG8zQAkiRiNIolMUcJEMdkDiYlFBy8+5xK86Hdxf56Np+SiBmP145tR
Ar8BhXHN6sNL0PGQI/9LirD68qotuyHZn/n5PvNPf0mD2NFAl4xKiKfrKJtLPEJ+
MhXrwL4q2f9c5UNS6fMf9ayarjwdltVGEARSJnlnWiVD6dubkX7eMcOSVLZbiEQV
/gw88rvv/EGQF8gsEt3jQpemGqsxKQLopd50rJ5MMKMFm/i9ZcMHkmAjXOa3SqJI
TZQ9z4XplHZucI2Vwxl0ZCyC36jrDGKNs///L58weazJL1FFKuF1pE7RzpMuGMiF
ScrFt1zi5FUlyOI7fd5qoTr3AriZrk8hBecSuI4GkEBws6BoIADZPGTYs32NvzmU
3p26VAXyE24+xKI4jx8cfx8MfBJ02sdM279Wd0nQmPGVVLLef4X80h5tSvfFqIgr
3g+7uwPtIzVowj0+V3lwEdCuYDUF4RBbSKJlrSTbBOZsFO3/NzE0bNNXzF+KY6k0
UuT5asKtiupg8JbKnupvbAG81vPELDInaOXUOip83w+Q7j9jy7MChCxKJQBxtx/B
7z0Z4vHVyFTq0te7pFyj9AmUd2aF1YGveMTS0q1AoUB+ayr8u9nO3MNvCTuX0LEG
VVoZ1y0nwd1S/kXCyGECyQtQ+BxIRNJ8aZLF9CCx90rypWLUHhkuMHTi3pmbsCzD
AUgNzlY1ZqRjDlVrgXXoLYH1OQMGEDuk03SlGufQ3KvPrEtSXM1xVMsdZhJ4e3JJ
Yf8L9CaMavzQ+UdM5SDyW6aSeFQ+Z4uCJ14s5xvIFtMGD39O+x+Z3bM9OCngP4AI
L/m4FmFFRABMA2SrBPmk3laDXwLkex5NvA3DCNPpc2Vi8bgR+ngbTDnej6Angj4Y
3aDVpBhZgR5sSYMFPLiF/CNeYMVz0kQzsZCZ0Zn8Nt1fky+o7J2oUcKI3vyhKfLc
G4pqgQoKc8S3Gh+3XEUeSO+ZB1tfQ/wVtWEjAjVUoZIAqKbNNPH7yHYhp7ApiiI0
57fuWA4FPF+oMjO0zZiucMs8/0CUPbCZgD8uceK6jzXuLGziVLFVpxpu1qQB3myT
Mw+c03Pk0BXcXcmVaHbomUdY4QsBGz+3i+ZobNbLLufS/q59K2+IcLyRy3qDUN3B
lOA9JByfV6rAXxdaIprx39ODaP7IkoZ0CSzlkmv5zJhjb8uuGu5uVHIFO9LY2Hb8
h9cUlarnRBGMCfzhUofc92vEz6kSi1SgveE3ZQXSUajDJp4a75bzqSIGciEH/onM
edKLx2gUsRAf/B+keEXRyq9DfBfcUY7Sd5qGVtYcYUxq/TlgMnQXow46xyg2+OLV
FaJPbLV5tUCAK8/KvYQW8D9K5A22mb5eLlYqmdNSRNN6XeVc4hr65fK04QdZVTch
qGFKIzuQXOdKG4oSF2GuIX0pdA1f1PWhQilrJpoC338/VZkCEkmaax5+KAVDO16e
UMSr5AOlFFnAojWUZxtWZCr8KKhJUcT6RiZsEcEZ43EcXVxAA6odTC+zJvsAU3d/
0+DYHCTHeNijPjkHkwugZ6Ed/0GMmy0CO01YONav1sEv2lDHVb8xUP+jM4G5BZz5
oVe0wmOZrgQPKb/On5UVoHVYzVGe3FKC5q6u6gu9KsZKv1APi6pWpQO5xV4i2mhb
pHbCAV1z19imSL+8gaX4GHNrsukc9Fd6K0/DudsslZI3pLqyDNkP7RZJjqU7DTez
fJM25/kAawn7tO9+OKGGVPLslJD5hEBa0BcFpVgCMetbLuD7+jpZ5MUH4afUbFQG
H3p8fMY9bOSN5W98hbp69xP0uf+wZj8494ac5L/vN+CcU10S3qiVcI5wIi8kjxFB
6v43edjrA3nPdmvLC1c3FjtoNhBFycXgRmNychh0Ibwrw2Mi5PQZhNyhADbeDSaR
8gb1Lt0cSSGZppttQw5l+FLIDoedvoO9zTHN1b8zyHW/8pwb9w3+p562qONXuUuL
Zxmi8SGLAzo0wmCX4SYopCTiBrMA02aeFw03TMufeAkXdgiwYgsCaHYdahF+9cGe
96Lxfm3DeYIidmTjRiBVtdk2znaCwLxTlaBjcOtXKPVu1M1iZRW0p/duLrGSsxQr
Hdx90TN/hIJ/w43jzo249sSqTLd/ON9r6YSLnBdWqZeReh/+nNeXNH9zAhUgFXkF
hxXAgCn/2A29uWi+6OCExO8sA42ARXte9JDkR+kDVXhC2xJim56E18Y/qmytYEGE
UEVzfUpBTBqjuYRxH5RxthhEBpUouS8S+ci9X7cOi3K1oUrMQu5ZkeBIHjASyfa8
4GDPtiLd/Cakgrhvne2HfkCo6BGKBuAfFJQTChLevf9LCSdLA13j0Xo+DiSCy+dB
57WIQTi5YPSq6SPLakxTrJdv+baCHji7MGoqJi5v5/hNboVHbmdnVnbzXHapCuvP
dC03G/UHvMNaaF37ervsF4IAYDaNQu2lvaChrtHV/FS/jIYemmUJ5A5m5UgQPxBP
JQIdhykLhGhgJaeGorqMhcfSSl6u7scCq1i9espP07focuOXiTI3l9nsFrLyaR/L
SK/UARpTlUEmcaINkGOUtAeF6fVYkcDrYcaboScTA8Nw1s0b7FF/0Pke9Sw6pu05
n4mc2ayTnKbrpTYADhRhDJnpiPZCvi7xiKiAmBrQxhkuBwu/Md86Jjs78VauKukY
odobJXhzep13ERRdd75URMsGJAT8vjq5jqGkv1PuikLQsu/9wIxyiphMSBZPhdSg
OrSB+CnYdX7Hwj/Uo1m1HKuijmkIj48eyRCbuYtzUEB5Q1B8A00VPyUa+ZmzES1X
pwCowmvF8uL+qzifUokDkjJ+vVpH3gcL5AOVZJS69ozHegxNhnaObJhZYETmMZ16
dHEtBit+ZfZC2Na/HVwtRrVReIsMM8GohSELLJATyrcBtKIhhKFetXmyg/HEOoWx
xQBcIdmmc2oqTEPO9GgiJjAabZgtbxoNJv7KsuwC48n1XojJW/mYS9E3DXm6u52X
Y7ca/xU0c2C420w7aA3oGGgv+zR8OPtKVSh0G+uWwrZbwlnT8OgTktPKoIvpAuwa
WtbwqpCr7udi1oPCdeOmqVFieOdd6zMJFEBRkdgobv/Qd39vsXhFWMC8kozVGEgJ
7FAxx5WPkjr/3IRyH+evZVi8ibN5bEmI51N8OvS7l3K2r5mny6RcY80+DoTKRQMv
0ys4w8OrsRfqxH5ETR4pE2RHEKji+NeyhRpaWSA1erDlQKRYm79JGNFYL4gDvId8
nNhTwuThNNeLsdNomYnxt3kY0SgtcIj+Rlmvn42wSAoqvjZ45qatY6AuZZ90/QwS
iy2Qp9RvGVnmJsV1VNaZQ4R6mrUxxvTQkuYoZIOTfUPHzlmpK6fabHcajBGCyEfT
qv72a2xjYqd510D92wHfK7zsOs5FsQJXlXn4KQvnopnzyjHvHmgDJUm64GRJVQXB
wrVLlclnghaZjZxTFI3NDrSix1Y4EYpDPeKYFPJ+5kXt/uO3tMK/0RZrmxzP5jwZ
P+ENIU3M/C7ZHuFtl1MrO3Ymgawsr998UJ3rHoXuq8YljJDYe50Nc6LfswpOBS/P
RIQG59+Qpsyp9JvrylaG40wKFtTx7tNPj7nt1G6EE5zK/sDpluIPmMG+mGhnxI1B
lIemORfyDBR0nXPgZugyc5BzXiSaTfdCKkI6wyW27z9+5mNjwqm3RKbt5CeokM0I
MqTNRIbmywtmOLENzx+dq7fe8ITDRvKMBAIuvJ1UHy8XfSorFQT/vVPnO/XHWlqq
5bc2X+Vzg3bPKXgunDqTXkZGcAdI8ibz5dTmzjQG5AFePBVlqDm8fvq02RvRnfDu
xWFVU1yco9vAx1g/iZvqb7EpGw8Bsu9a4ur2c2c4xWf3ZsZupZGNqE0DU9j4XVDQ
Pth++GA+pZwBSuZvvHvUPeZyb1zkii+C58WR8E8guCCJoStPHo0jLXctV1I7IFKC
LqgITiz1LJZyCisgJChaN36z1ADFGCpJoikwDabpdhDD9R0pR1EHY2YdSNHkhk5T
zkIF88Jv8xUWSikJTmams8HE7f41hKZc8+AR+sMiB2IcQttWrDGlf7CedaQnUqtz
E/CA2fGgYm47T/KREdREUvdyMEXDxV4OMl88w/tGrKIvZ9PO5UHmefnXfjprwxdB
wiFjoI+MY56VMWIO+H4bZhQfvLCIkOaNDfFww7YxBdMJVEr5eg8hjW5SpiNc8nNm
4p9mI+VzHm0b/VP0t6CGABC7oGsrbhceGvStBjuZysvZz/004Cu9xT/0V/vGD6w4
pWS0r9boEHlmVSrW5g9Zey7OqtHid2shcCR8yURpOARq++/ZxFIkA4MiQ08zFSgV
oELmFKzAe19SS2eWR76QmkM3ZKRfOqMjWwu6HBNJkSbn555F6C7+NAQ7Smh3V8qA
LP9VBqjCS+OhqC5r8T+4Ev2xNZz/WI2ejxARiGe7r0VCh9pJJSevUWPSRL2gdZEV
//SFAOdldsS4IcuEfNJu9XfUbU3BUFXEsGkmbMuYEG3Oq32z9l2VDiZpkrD3N1V3
0Egn7XtSzGFd128Io4mn+7anzusLfXZE4IR2lu+di0WICqF3tfuoRXbdLbnWTKC5
m1yaXFKm0gvs6LJn02ZmYIEwti/uRMTxHYBStY3cO2Ur2nqqBV38GVLb4rbzRtG+
gSiBv1KqRHnW8F+a9Vm6Dd2IDp0mohAjKIjzHnkdkxRNR0V5orki+LwYLEBZRHAm
+YxQWII20f/ap357BaVx/N6V/2i8XY4J40HoNxA9pHhyCbzZCQaurp9/t1NiOIYU
SVq1TmVpPJ2wWH3f9JM8hfbe8/2xJYaOgOjYrlJtx1/B9O9DjOXL1fvqN2+QVaJv
a3jgs+mkeIHpcLPtIaMiX4GjzTovmhDBzzm4pXIwzZPH9o7Xf602wv8kf9kS+1lP
JPBDhtGEg6w19MBcFHDKY6hfvTvU4JPsolZfpYlAsURYg//XYyrSwSL5BLe3B6tZ
pWSzd6uV0nCBHtDOik1AskZeaoK64hdTQqSWX/cD2Vc5JclejZ9t44e7cs0MPCUh
iaGWH7VILuBD5gyw/XIzIin/6NCW+XJ0UPuH8XxYSugS8BBRGrqJQf2YfZD/JVUc
jzYVT4JiORFxWDnnYF8xu+Yy0TAygoKS4oXaiH0kE2tH+73RIqU25fPVDcPIpL5y
4H6kmIIm4389CU1GFIwhUFY5PW4beEQvF8o4tiunIQdH+47D0+hptNUhaOFTlYMC
cjCD+vQGA9qeoO78EE3S1vdR4Sp3IHRgPhWViPm/aadcxN5QkmfujhtIiTk9D3eA
NjMnnQVTjMLVxO4klwbdMdctHkWEGUTVfS7jmLsARPDEERkjXXG8MwAHIcqwobYd
xgyF1n6rYtbrKy7YVYiC84QjStP4KSd1Z0QJFBDgS11FDLvzS3bzSaEVW2aDGjrP
jWhW2tiQMRXiGj9psjOQvfxOEI2IAklnQQPCNJJYknmxLtDdsMzhnsS7vTD5wGKw
n/jLTPWlOGF5esvk6skX94uMVxhcY1CmVPWrKZXh+ks+QjJ74Dk8oAKvXYjSfCCu
2bt4m97XGh6cEgkjHjadK2I0y+hmOzwfA9WO92fhzUIQKCtkP1Iw+RC9arQ0gYiQ
cnZFzYxk0oEP28wf7a7TvEYWv2cylynnv/grwe9xIaQryxCTMhAdPqkBX9zQzQv7
YJEXAFbL91qbb36HWnrNu3zjRAQAIpwCIoCMdsZxksj4fqLA4ZEJnNJsPQ20ia0I
2WPAbZDOid/c+07KiHGA4Srb7BIwMIv5nQg1GiB6GBaqx0Jo6vhWYnSgChZ6TKN5
fQpSsaV71paeePXwueSNHMEMy8dp3gbe/qED03jkrliQq0dok2OWnw7uujsV5v2P
pJhcyPf7A03JwgbfsHdvA3XGeRera7MKxPIYCvXqLLhFiP/svrhdGTtLFdVHdKLU
j8gZ95O9w1XLVSUPVQVmc8xSlvEviHSv+Pir4p/zaJ4B+BhAM7ouXWCGZlvhHpyT
hdHd2IFk57drcGnB4/eqnZMcl/DU8PvKPYVKYHoLt+AmYBEKTitB9J2AXwe69gC8
8ZnhyKpPr3Hiixi4A9/mFOOuXZp3cTksCu0DvoXFQxQ6CvEGHhidzPzjvX6iSnyj
72mLil1Lbf+/WWDAGm+n8EXcpfXCcvXxQo+yJXiaK9BiYfx0v1v22OAyP6yFggDF
EzW5gLaG22I976t+fOW9MBFvc9RXASgtHZKIPvcmHusoPoBWdN15rJKNfc9wME1m
q6fjOUDqOc1dg4AvPqwMnFZI1NvnoRdOa26gbSST4ermZvM9CRKtsjbkKpzFdiqM
H6dmtoEP1qRbGeK5j6l4tWTTELUx1Fcrp0zTggFIiyEiQEUOp0G39nnpRcMeBZBE
csoYT2ggzzUDDOVexbJq/H5ABgu5EKqqfXtm+ledDi9dA21zLfq0FkyQnfTly3aT
s+etV+zOXJrSnG5FktJRQVfwqJaroyEdqyXfj+RRej5nZZYD5n2UDNrkZ0neEMXL
iICIeJ3oxCv/BmRscDUMrQpJTHHLxstyqYYZXzGtzA20yAErvuxzhJ53JtXktlDg
S/mPRPmlHxp6CCJiAh0rPpxOJOsQFtObdc1DnRFXLwc5YR09/4y/IsDpsfgbhoiX
3mDX5bcKiVSISR5AqL0TOi8o8JSEy8XBYBXBjRoBl5bp7Py43ByWU8osXroR9MmK
31sPkHkfoW0BZdVcmiqthhIDaJpMsw1pdF/q3xj0AbpsWy8t365esDQhMYcH8Ygc
vIBOKUPtsWfEV9gs0qyMy2hGivuxlP5jK1flwVT+JC1LbEjArPHE1KsJ2NaWhfrs
/TDQu0KxyPWyNXIMtc9AxvQd1HyLnA4XVJanU/rkh/G40jNlXPbbLw66xRiXNXsG
rRDTlmVToOBaStGoTRStCmBF1iXjubpVmIN4zS4sporDx8OEZfcE3dhuWOYJkl3a
K+vkG5Vc5OpYgNgxMQz6xmfGtuFGBJoceQ6SX1E2n8VlAcZwdjQ+/wyMF7Ju4/y4
DRlr8rStsb0evK7Ic8TZzPBplxTWZpkSSiw+VoyIiB/wBmA7QidzISGJ/sosZMLz
xkWMwmb9hHRK+pqS2TyGJSx4lCYG50bqHBdidm9CYww0XHbvZtoO3PL0SC8IB1Jq
B3l2zrGERPzxHYTVhVJOmTxuYuIHti+QZFIuhIXIOzn2b3OmBQ8o3JbKMC5GtgAb
den1LGQrI0XTpKC1UFSSX2uKh1t8m783ZhVuSfnOdoLFhUDJnypEQgsHlMdNvS3j
irg1txNi0ErrjZZzSTWZfP+WlzgCnMRzdHnIcntEGTEAKhtPVJv1NPLV2lS88zI1
/GlkW9KpyXAR87ASujksZ622wlEiw6T7fwnzA8Ba/MNBycmTS9FO4gZ6rFGnV+Wb
Z9xhqonsGDW7/UMmcIqo8PEO0ttIACVz400qXx7wrN5l68kODz4KvS1S3shOsk89
/NbeoJ/JIM/t65PBfSoP+PU9NMP+bOe3JQOnDYfQ3fCIybN3T6JcbIc7OQ0PYy3u
dsZMSfhxv6hoZssVpQjTa8NuHimFZpewIs10/TxCOvWPw6zay0FBH2s1T4KH/SS9
/5FW47C4SMMNyR6aaHud+NV6z3/Xmx0l9rKSOwGx0KGfmo4TLuY34yNnZE5XZ6WQ
+G1/VuBrYIdYxsvO+eJJEAi/yjxxS3h05TsF1JBakCM9GAdLUMPmS1xoOEGRKBOA
gLwyQre4inlJCpHGB8+/HzIS9aQ6puThEtFXRNWnzZpKj7NZwKbZASCQNjHNJhgI
X6A2qEg1l58GtHoXF+3PJwmxl2Hu+u6e+0/m1e4hjFkUav33zLsjdUNF6w8KN92S
jQVs6mn++1A7hmlBlRwDQlZ/o//p+QDeu+M6JkTBFes4c9/JnABXX6msyIiIl2S3
/sh4mrdTldXuUCoTV3RCwsHHOnHiBHyB7nX9KmUJycf+h1T0zyQ6NJcxWcSsBRFY
UKv8LxzNpYY2HuVO4aXuOyTOKP4CzzJPT9skdH15DGQ0X0yObILPCwl+qfYdE3Ex
wQPqFVXNKXSPzny4C0njWvKvtUfqWdQVKLM0eXr9nYpoKDkj1huHwoj9NCEWiiiB
eRFZx8crDE84sqDO1+eSS7DPLevxt9NioPAEQyR4bv7A3iECjEPVuZyN+sgLVjvX
vJEsmV0c/v+K4SoNKVI78mgSiIBte5OFfHpxHpuoYwiDUU2lr8Nca4ut47Q9dbYT
5wN2Vwv65YiC8C989p/xwaOAR4PM9oeCGSFVLH+tevBgDemBH+7Dqx194w14cYEU
ww4BGcrw5PNyw+9S2wszTTqr6D1L25ZpBI3IGltDHYsNqBvP6rs3cvLEZcd4mm+M
X5lyiQBMCNdu15AVnVnGCE01gVI6Ak3JRsW+jFlfUckScBVOaksRS8U3JqG+Kb1G
HLZb2ydSIVlY9Is2EFY3159QJZFQmDWqgE00iISRP6e8T/q7u6nYL1h2CkoEMylH
zPx1vKPoLzuz/0heozf1w7Nc766KZ1T7v+JhXPwbZAPHd1af0j3Ezign+faYoG9N
JjTLebeUzV3Y1cyI5TnAQeDK2vXrpVXj36TIJSDAR0IXnc6JUcGwOmvsecckvom8
TN0uc9uTNq19LEIrS5V5iNyft7e6DR5flZdkaPBQytynUoRd3VbG1yiKG3UO9yhH
7XEoVhBJXfefcHPnah2ZjDzLnaMU28ERee2vflcYk16e4e3elB+FRMVlp2Ao+GkI
liF/vm9VMZJEjQ7wMW0BxFcAdhlOs7uka+8sthDQor3zSTt1Xq05XFhYUA7CWBVe
pSMEn10CXheoHPVUKq469hMr9M2OYkzAxNFpHJ7ktjVu1OimODOK1fdop8CLdMeJ
SDVjd4hQRw+6sWdXEk00dKPOdn4B4z1BuGyXx/TZACc2gDFwjP2jNUZhPlqXu3uX
U1/1Pw/qqFaj2AcxhQhDbt0nVXyF4c8xQ9fLgsXajFdoRzLOeHrAjPt+7bFN93tR
hWZG3KM9LlhYZsufrLCppJvBDFhGLB7kNnbgba0NR7soafTlmW2RHtFi0ArrxUA2
eo9OJi6KHcYatn48dLq1btKnT5QNo5k36cqdclkIroJjoMOkp9MLP7gF9M4e98YK
Mxp2ErTr6VB84c0yZbXfXzWA1t4CJmRh4redtlSaGXy866ksMMByDTmG4BXN38FF
GxDRCYp1sahLE8eIT0IASdIU1s6+StTFe3xSjBTY7q2HET6ziCzpe7ha/yJ4zrdD
/gxOAojYbJ/p6M0Mz2hxx1U1/DVB/Up3e+3tMyMhbeLElv7yB+nfgISHmrU74Fcv
EO4qLP6ofjp7YZrU386//GALrFG/Hsu1vV5PrtJUggor1G8txfX+Vt4yXJD4PSqc
F5yrdshXoropvQ4UW6+rQxmPbQfUmKRNiYaBstgr9nA6sf3BuWfXFyD9iT/p8plX
Ke2PxWMMZzah9bgLFg9HOUTeQTFKZ66ZUDUUMHV3fx/hnp/qWpF2rhfpDqXQ7pAx
T9KeNB1D5+6u3LcR7e/Cmlstb+LdBSbp6MY1yL5wAwYzwwJ/O0/HTgb9SUC7Z1KT
5XvHVw6lcxLYKI3zs1rlRsI4at8xyBCVBx+GPATcWrSO/xCNr9jjTNpsbg3Vc3MP
pFLAZ8uZ25qfqWdFKftWV8J4/eoBGxgee1OEpiIGyleJAx+nQ0pCE0VYTT2XkvN3
rud3zY0fnBa87Ozv0JFvIviZBgSRnSQrm59SfzpKoK1i2mQrDu7JvWSAYUm30kOJ
aafd/+N6Y4hqTDdEVr9DuP7iT41nXfjiM41EWyjL6gHTWlMJJEXR//ToMVM1hRB3
RF9QxEys7kfJZsB0B3L7TFIhpD407H34K+jMg9vtkshFCUrSFRKoe2HjbrZh9xNh
xNLxLbgWVcvXUMpLpDgdIAJU0BLqq1goc36WGwUoIhSzr04FIUyxc3qc1hSkgkHR
YNI63tM00BAjBJEwQZBM7ND5IGAE2Bv54kqiJv6aVXUVCZd/AXGtXQcWQUrJ7Mfb
Z1TULY4C0gKiOSBRGuM/q4vS/8NCk34UVc1AXalTVr3oBxgbAxsa9Gnlmbuk2Ha2
hz6N881e/xdzPM2768TaV4h/wfjlvBsXVFZb3xKd9lzMTJcVAhhfYLZSbLxjL5jp
/U5idqu/Tb1XgKc4+QtwDltJJ9fiRxcuGbqnK79upFMNUH8eIiMAjYBfAiAVvhpl
swBSPKApfVwD0ybDqxXa6TLVaBbk5RQsQZwV26rZDGO6IUh/hys2okF22lQVMRqY
MpbggrJzuowXqqP8pbq7v4fOUs04Z2/9DOC9xr2R5bUnVtH4fPqCYQQ5I6pjO0jL
ywyJW84qGVqLTbHyzV0kc5lMkG6GBvuteu2tOtdFj8wceZ9/3RHehInxJteg3eDv
VNFeCHARSFi7b196H1Lzl5rdJZ/37PgmJFgrozH97WoNKskS4+B9p4CT/qduFgdm
L5IRnq7EI0XvsSRwNxo2qS9HEWFyGBwmIUSTbzTqS7oz48SbsVzB/3EJOHw8/CGa
xwp+Da6htT0jN27+lwgpK/uBEFXIBLZX5u/YoCyhuHX+au5vnteQX/R6yurB9Ekb
yijpR/VhXt4Lw1xTqd/dV0yD5QbLqq9pDchpvNi+WnhR8ylsOecnfq1mzsy20qcL
Zsp453wkxpnuhQC04Lnu7FKALbEYQ9AspRzdTTPJWzLomIeWxb+5AsXe05+YIQOb
laDR133S3b7IAe4/iwb1AehGL4DY5J0YhPPM9XCcGno+8TSiW0ENMcNMJewqvDhY
IuKgs6zY3Yqi6fdKAiumbRgrl/l1C/p4IgBu/iTNhplYG57dsmxSeV2fnrg5T+9N
OwkgYMf/Kb6i/thP58fQw1HS0gjm/ZRAxiLWN6M3xigwBRePKYSNf3Rbo/QbxM80
5oSOevA3V7EGo83PseeHAh4pi/908NPfxFSQPeY1jrLlUGVdouvl1kIsseNiXIIH
TZQnq+CHCCToYp62//m21bx11YufCRgIIHhng9I1BLxgwlzNcP8PGdYShlqcMIlE
AmXMCnelWxl88VCM6SuDbMP4c4lugCfHzPX5Pie+QHj3yW8qK/s8a5FtEXbjYImQ
9zsp/leXs/sPFRICx1Zs2ULHsMCNeR/EosKSr1NSTf/Of/hWT/j1KrcPCfxtfEbs
Ngs4rfLP/lMZnWgsOAPrBAM8CS+xtkt6f/q1ksbU68Fn9psah1T72Cghpl6njmKn
ASL2lobAFYX87RDr8TOSdHXZyHxe4u/r2+793VS04Q0340CSeFp3oW6jKdjw6ZwR
2TO4uULgBpR0PXvkxLmW0Aa/rKanenBybYvUvY9tyP+YwBCqRjvIrbrR49VaGsYb
QilsKu0/6xtaFF/UjVGFsplehPFFh5wmceWvD40QPk9SM40qB+R9vb8zThdOc4y3
r3+qSotoAleAPuB/GgrY6xBmyQu1D+LgZElVU5nak7Jnoz9z2TCFyqy4jo/OI59H
XUec/WZ6ASxyWAHPkVYeMlXAD19rRWI2FUNNOwn7PIXNWV7iK+S2XAosQHPQtHJ9
KUYJX+rRzNElCKKkkjsqIcrAcgBhEhP2ZE1x4pqoLgrk3h5xMEeZbrLt6CdMtrx5
sIOKy57tswHCHotS8YRRtAa55uURox8Q1WtAcmihvrkqXhk3XBwY/mgXTLtLr6hy
R8y2Qt/39QnT9HzN1pnSioHdf+0MvycqGHjmFLQxv9Ma6/lWPEWygTYd82LvsJ+K
1rHBSDOMn4GeTOUYv/rW4SpG7j1KdQtXtjGpLA+Kkr+rh2F0kJqOxMefahZ2dVKA
ykqs54yt9ekdRoVi76SWazUNxABL9HvbWt72u/Uchh66WwoejW0McyaoA5QSYsr8
bC+qS1XrGXXbhgFlr7bRyiV1z0xVr2xcbb9WLUelgl5X5Zy8sBbVVXFm1pAgb00L
j6JJqSxO/4eDGBgFYGLok5MDJyr3U5v7U8CORZlF5HLnwXg7tEZSeyDJbqWryIqy
ZXW+BWffsK80lxTZTYQ76yVUpFyU+tg/YXYU4HaNJJjjKdtRh0smeGSPFke797G5
V3fOg6BabRFqLIbEzTj1g++GmcwgOcZzt7gzF2gEc5mI/L6UddyrSf5PiNuaLLKg
3HghrySs4KKfWDRyWvoXEBVxwlyD0/e4ioLwHbhbF0TUtoNdnESi3HtKQCEGVeNQ
2cES+VHC9Wn4xSuZ2IffQUIwtuZC78qzSN6DFV6n+LwsLdIRXL/ZcJZAjDBrD4aK
tKKvnlEOtTX+zgnAiAWJn0U6Uy2jjBxV82AkF7adiYD9KfFZSq8rBkRSh0eIDvHz
o97F/gNWty2lGrtYO0+3EyyZJdHw0N7Gv9eCiONO+iHXDL+6ScaH8kAY/rf0PWCV
sfv/pNxrc4uK+zzz9zuaGXojYKYPoRePE9hC67VmczXEicTLVnPo7LuG7+Ns/dLC
c7MvhkS60h2QjpVOXlzjXs3s81n4cWt55XAp6Nu1e1C/KnG3ggceAWDFCM+Imnp3
yZMIGO1dA4LrYOZSa0WFR/rqy3EP2jfsvUkVE+xHa8T+QOEOdV26OyHhgBTSos7K
3mv3drAp/pu2cxzD3QaEy3jlHbKqkX60eLW2vLPgH8jnPnWnmQDhYnTvyrLq1LVo
Jgl2t642qHH6PoeJIdcXZoJnYkdA1arYfTI+53p2PbNGK50DBzFfje9hVHEc4riA
RV7XDifTGXTyccXRBeuN1jf/g9qBkEz0qFisjpdzXNmn2pih/WWwhLJ2OOqbMnEX
cD6ic0OdV1QhIJLG+luXMHSWA+gLUVCyQyb0ylYqqbrvWPHyxJPBGqFZCUqgHlSq
Z1sdEwdHO3DPbiKod87g7X2SfKgyHY8WhYqWAZKnlpkl7M2lsu4TQqtqZ/uvRRIJ
S7QisWOIvukZkCLE/QKz3UcIbXuW7jxlnQpw0FML/Wk0N0E5bxms9GZXkn/PIdev
8aYZGK1koGO702f3qAirE8lQesaHoIDw0u5S85KRZPyFi8sYXVXzI//UlLJuQkKj
ULhxjb6dojU+W1Cp7hYwQmbzXCSBtl2KGx0mB0n/fyGaAbhgHjCUcXvA1L+zHbMx
H3oHHVS8aikXrc9mK0c5/sC0jX+BRR08O42Q/uhMNCf3x4+NZOdEC8eQW3zqmMn1
DNvwEOHmtHR0LRRpYx+0fFfyINMmT0s5DimHrC+qnJ+45xQgixWzFw12UJR9CLFr
X9vPLmigY+q3Ijtc92FeMGhkNdfDLlio+wBbgwODgb9/twUe4c422amPOd+jxUGP
WXFWLaVx38z+GkmC7YhN7RRpm/vkgMJMtggZ3H/wyBZrQjiZIuCjMAFH5kATy21P
Yz3fViBXmH2C4BPT2ZBnyPam6RIYLjMWBcZFpDWodXsN5VJfA8wvYp0+DLo1aNfI
LzjLNsF7k8XrfIjRLX2NcbhbpTrdnn1/5IXsxT+RT7Na4aG8Zy7V5ZgqzvmGN3Fx
NSW4R1cvbryn5A5BNGJtO+E4OL1kyG6wxL5ILa1mdhAJv6E3/UieJBrpBe47GE1E
Wqboz8Iq4uIFli5q0Hkrzxx0F4+YM//zy3/Uoyuqec1uGm6umGG6HQugytahAS7w
D5kd/AZ3VztDUTOHVCj468H2EVrONaPY0itYfM/gI+GJZ2WMcPPDRAl5ePArjRC8
gaaJhp47F2cv2TaC84SEQu+Oaln1SuLtD8vgEMWKixOHHwRHI4V2EUvR9QxXlO8s
AQ2eS8uA0tPBRAXitTal9QsUa3+kV3bXphnAVhEoYnSvv6CR9hSxe3aLp/N/D9ZQ
v8F0bwown7c/mBvbDwymcJnxf9hPouOYU6cjtRFM/Q8mYvVb53FDHpguS6joCFCc
klsr8/Nx+8OiV2NhX1gcAuLT536raLOGzPxYQE0XW1fO9A/EEmyCDC2ZmRA/HwOp
h9oThSZh4TMQiMwK27SyVbnBYqRNDP0Oe18IFUw+w2SAWKQOEL6qYyYxIYuTZUtI
mlqEsTuHXO2f3zqtlV7PML1m+FjLaIXEDOZVp06FdgsPrKhjZ2yoQ/JsWgNFnJbC
Ww9JJQjkdD46sMpKVq6WzltO5kfJd5f6whVk+hx6809/0S85npAGkCcvMIItjqqB
KhIevDvzhlU9KT1xv/ithWplmQQxCms8wHBnFX4SyiXEqliuwS4Bt/YNFNHXW8m1
AYZxOo1bylBtELGIcQEvo3gSmTSthGMLKLfR7sh+Auo8N2pv0iuUj58hO3tYhtk3
O8JFCUnL1h9HUePc5uSwGhkGYaHIWT4o1Uz3Z938oAbDzWm5gqNGT74kz5nONso2
X7ULJs/gnT88wWdBomYox79DsSG8zrxyseP37huaMfBa0jbv/6BCybgTcnSoP+b/
BB/9KoZvarXiQRM3sU0Cy/csahakbW5QH0DGwyyr/5qfpFKqSnWCZf+eOvbJbr47
sxXwxj5LY7iUGwiVI8jYhW4RqN9wi9AAzr7ni2QJVwkb3z9I5WOhcYUO2zFVR7D1
Ib1Kr64PWZ3lCqtJsHU27zVn0gS/yYdOlsxtKFEjLmyozioSrSsZRGH11s5Q42Vi
kMUcbmIK2VsvS3uUpU2n6jqfVgvxvahTWwLL+VbfyDtMsd7zAVWRx1HCURr2ik7e
2pJwq29e7FFvAb2VboXw4gqEI65HUSqdp44wXKDYfOgFbd2RE4H105QC9BzxMOid
klRbb6LRRs5TBJkhpwzfxjMA1OKcoWOEJ0vtTwZkntoUifu125+u4bh1dbHxkxox
7CoFv6ZKeEXMH2H2ImP1O1HuBLXJ+280di/BpS8mhJwrZ44BKoy0TTSYjJcDTQlr
sZ8tNYVocrRLRL8YEJ+9s4+mJmfFlH67tHNvZTwnAkPaPzJeu1k9/y8w9jHSSRDT
DSATYdE6ttVH7k5jsX098poTmo+HA65o6+m8TB+Xqhtjyj93qGKG75KL9/AdGry3
QX3JP+WJDhG3Wy3929qRRqO43fmeBTcvUz84P/I1K97dSZQcd0B/3F6XbjTXgMGB
mUwV3RZN+o4iJIA0zDksnR3+6xN9a9FrZuPEsRDVJeAtaeoC4oV/Cc6hMCMk+6nW
zk+mGGbSqJYjKXhjOR5R49x/zVeX9QHBz3d6KSYlq9xkftio2Pqip0zGxnURdbVm
2JPRk6q2aeAF/g+gEMWTony9/0VlKKn3FXPLH727EmAxqDCVdGm8ugIioguqH8BF
d4e4fjKDoRTdgmHS55OEHvXuWerLeOgZTWp41tYEreIdWf8MdlZJb7+EFamAw60U
gn9nAISsSDPuz5TavdIF/qtOjFLUttnBY2gJ5FuTSPVGFwdiKK0yIxNezvywe9X0
6psVWIfpi85y9YnRiTeH3tKi2oFPwJG72VX4Hdjg4K1VjhpUN5WRbVbYk/d2wadX
dRIl11t7kBaJmQpMR9nSjxLOfUpsNja9QGKbH+L8akRfNOWj001oBt4QfPIQH/Vi
efYCWmKKTBCYDeqLVzDIKCBcRbXNLqA6BqSOpN102KMbF2PEDuMXDLzvGYy9ktz/
njBJ7jsB/7Ir3SnBj2GlnM3tzIL8ACKc8Irwd29YK9mciIA9IcXZPBIXOVYCY/Uk
ykPeCli7SzWH3yx0B3OvyY0y6lrZt2xvR+ymf35nuJ96otEshXNWiIhNsuAuZmdU
k8kEPbQ9PtcBFwHYchb7JnngkVj78UN0Toz4eJn2osQYygtIWvPMJlSVfcqHcw7b
cOAUHwwhIf7lmkCGtQgZCNPv2Dt6jkL1r3ZC35RuRavUkK7AoRwDatYxlxKzZG1x
BPbMWQBs/QZQu7lG830akhbxQwpISuYyzuqSzK/p/+GklYj9UvUmBUuxrvnr76zL
7jvleSHifuQOEzKbXX0RqXwfLuIo9IFXYpl8KLqzaWLsCqqDFGpBKZl9EFLcR+bn
vzFyJ8cGj3FQ8tSjrenvqWPTlahoT09A9puE7VndhQPrNAbfnJzwBMzgYmxxUlzv
xK7ws4clXk4faZdnSnVjiR90J7whpIh8Y4Tdgk+khiGmzmlMExVNnkiNsyNjYMpp
Sc1muGvrKOAz5uoFNVpxBiUQbKmpV8LqdtRRafzUM5yyxdt6QRKl/dscC7OsIZ38
qF2T2YX4ZnssTKhM3qHetk4X/Wf6IeF8TDQmOkM3rWr2VF5vj7optQx2s/gdnHDH
mPRpT9eWRISh9jz+1OavRVfWQwLpwWSzcwMb/oP4oAd8CVnhEZHyrCEphFw49c6d
1RNCYYtnP6pxaIGkvAQvE9WXpjU0BjXhk3S4ZZXm7tDhTGswMo8BHUZh9NZPXNVe
QUR6T7LtddavZ65oTPj8C+buIdBfSkC1yemnZks59wHN+9WWQg1wV9xxxCZeAMd1
Ak45wFoqOUNbbBAbZYj9IMO7XEHV5fRIffGgU19pQVKn6FI5BpYbZ2Kqga89lQCO
n1bsOUldCfIIWbXBviFyThLukZ9zeN/ZJSfXdg41a9uDJod3Q/Wls0dwb1lEMXJ8
RjmBm9AIAgAZ4VhLg3fI3cOHHYxAAfPJ0Hkasqh8xTHov2h7QSl2JA9164NF6I65
B04EF1YGKf/vEKppdKFhLatYXnoJTclc5PdYBGwaItVyCMxAd/P1jG8oNW+ZRV/u
jjNz7ufTvPUw098NplNr818PoXHhb5Olr4L1I78KMG+bS7xCFNGO9CDnZkqy5djM
8JNem+eE+VYC6atMk3zHSeAFGM9f2GZVrkHpBHJ+/LrKkvKl3TePqJHfX+IoIVqV
T6wA5QFYMNmw02BhpKHAGc2pxeAtrW+p8IpsOksoUfgC1xPMDzPXi8OofOFNXl5r
uHYIna01+rtbx/4pZlYKMlLyC9rI7SpHULu1bZHBLdHkaj14UL6n0ZV+FCBlorbM
WN9f1INkDJC77zzfsG6zjCtYe+zFSfferNUtYEpCb7uxOlkpBq48Vu9D1HlXUNU3
0qoFFX42omsig6bijo7Ru0de1PGFsn+8Col5zZ1GhgZMovOlXFIlF0fPcGgU1ZqC
i961UI6YWDC7u84FxBLjbBUfjaXJukqh6WTbgfTEmFs699WxQRQoIcm9/DdWPDc1
6qRox7GOyRC+wmRLTMhSwkaHrCdx4JHVryAqmv68nXhMzgRCxKW8orXrfEn9IuYC
DP04cgDHaYogt9QrwMZ+W0HkcUlYqegBN6b7TxZ/Ki2fE98frPhvLdWd6kh5RfQC
LIwco7/jyJ1PMn4u9OOvQ1q8juBtl6HnaOyLHlgAHr3CAYvAfLuiCcMxV15wmscJ
3zk4eHMDHi0YxM7SBSo2FiLzVPMieFUMDBbnfgBfB7Cupg4QIYrb2k4lMzSciisZ
kH4WbuzxTmidbSC7RDKhsca6Ocw0Wsx9q7fLG6xtRSCrJbdpkDXE1els1EyxsTfZ
da6LQ8qK8bA6EZS629GzcbrxPj2LKIYOvTX2ToF0j5/AeOZ9J5R2bE+6UDeSw36V
Q4F28ii2r7BMniaWTGx0vBCTPBil7cCtrbzYCerstAdcHY4H8RPsvm/Alw+RGLtc
HOqePzzJjmpShpp3UgV57twSiueJuRsfx4EOjwlcNH6yt40CsnOuarFBq+ThdjFM
UHFbjj4PXs0uvEE//0BsSAIQRRmQBmxSgHOaaKxTdP01RH6cFuCph/d7k+N3aJs1
ve4oq0rprVgYbP8KXFc1wWVJVyrVjkBo1jZlpxX+u7UtVH/gh/+Q0YoHvUeYgvO+
+kt+k4zOL7zTug6gtEBelRhbEvgacMvOi1zoBTRNcOWkgfOhwyVN2XybRqrTxSqV
E/HOHEuqYKMH4bGj1KXtNbMVT8nH+rY3Zmg7BJIi3Q5tbwYqquQqj/IDYa0jbdI2
QXA/o7f3v9DSnddFeEar9RbNCvrN9az51ASScuSR9McE0DB26ZQrYDORgut9wV46
P9cVoDIEuzrcSm+Wv1wOyNiDO5O827XDI0Yhw0T89BzhENnoF4GUv9otJLv5ggVO
oyysh7orrehubTiI7rKY8GMfKeu+j3jwrnwiABFen3169562WHu+DW1IWsax4NWS
XpIi0/W8KfM6aRxir4O+JrltKb5v7NJ/XOEULJWuitPICz5ZrYD46YDAY11UNHhA
YTryTDNgcmCBCXg4ciLd4ifDIJ5xWtxk3XAlSSLVUP8N9pwLolGn6VdTpYSDK95j
WUOjqfLHIrJCAqi6FM7v4/XfcPA2+UwUQm+TZQeYBl3/YO8CzybDrJA9y4DptsdM
pUE2lbMIHk/5AAF5RWxDBR2SO7HXdjBBELxI8MqWtonB9+ExHAx1u5sJl5U3Ay3x
DioF2Izool992sfVyRqXOnvBVICUsE4e0DfVjXZplr/yCv9gkgl0DjFCqLg/dge1
/GcOqx24teyCslAp9p1absXif88jKtWPZ8t7A4BMaWR/1qPH7HdMIp/8nxa5++eW
yBrfK+qyDaCkIU0bnCqx9j5B+2cjLq2g/bMgKFpV+j1kH0FqugC/x8wH92MCygzs
TNjrsDoxpuY//wV+UrkoCRB8irJtLMnugG+bTadn+pIRFlVrY9zZkhnn4m7hnmm6
lc85wGNmfGbe1HILfb7yt8wPVMYhrA8ovKlsMJivKTmbDsFQ9wfSjii/HL01+I55
nvMRIRiJ6r1zVpB4z42UpsRnPWO3RCbdConQonROTPMbLJhejuI3zPEBa/1xpCcV
98EsqwmoIJe24lCEiSBXNLei8cB89C423kUTTYGdfRQVtREqQ0y3b3OUUB5ZFiNE
BNIevJXSfovIMG822FhtWlgVmPsXWsTK0//ICPfnmk1kDPc6Pt1aFJoDXgQclNz5
Qt8jEbWH6Yxme3KQtsXKWYus4VeIoZBHOTOGTZSt4hVb75+bMPYoLNxSyyJyrWyR
R0QGVg2BOC9sGJjf8dOG2hXj8rxpNd2SJqX8A3kpxbtbsInNNePVvYyv7FuXzUD6
d7IB99znilXGRkwwa0GTIZZEdDrWF8yUhifQP/ol/FMDKFjAN4L+WXalcBRQv/fi
LJE5jkv7SEnn7YXslZiE3OdiberOEqnqhBKAGWJiEyYHQ2ufR/5AXaYunYAhC5Ar
MJi+ylr7iV2c4yd+GmfyrHHWxquCL3VAWohkUYkV1ubg2amK/LdkhRm8AW67npaT
2Pwp0QCrcQ4eq9rVKeftjMlBxsJQpAtXtiV97b580Ro3WXqoOzQ4u0s2yRBUcnxN
b+bqpBr4GrujvHNGjcNY++P8sM9ZnPnIj5ZXfj/iorgYN0SIT8B5LP0bTwMsMq6F
oNKHKKUjJL9ZlZQWmYd4wVxfCa72G5jcjjKGR1j64rQTCiSyBw+ypT52Pbkv7IP9
eLQ120PKtP83RyUMgMQQp+e1uLmf4DKOuCpxThF7MiIfnfNePVMUxUSqVzd5trbk
LxdQFRGQL7y0AU+aiFJl8nSbXIxWla4yA88eDQRbJJGlYQsVYW0Ptk3anvDSn/kH
meJiBf+R/DtbRmwGQdSj//9fLjRYRSK2Pq5xjx16gssdlRtwQsBD9OGxjoA3jPw5
TGzk/z8KZWqe/EIZoKz2adfp4rmL/opuPbXhsc8JtsApF13vMNt7SiXYCRXH9uhJ
3znPCi1lTcaiGUl0KtyXpZ8CEdnkZrQh8dgmBidQAoXPAIsqq8tN112coOoqgAbK
+Bo4hRfKPcZxP6arqDE77KqtQlUVlSvz4sn3tKDQmXJarDBJdJ2qLGlKDBNxKO1y
HwPU+khm63Kfpfjs4QW+0Sp9Y/iy+JE9Aw6ob5ePcBiv3eZc/vMPtsVxKQePYnrz
QSkqW9Y8wBi8sz/l8wN36/UJh7kZBOa8VfA4Xkesv3s5NuvNMPKN+MMO1EPbS1HL
H/x8qK2goTGDI06GNzGO47T/X6xl1uj+thtWIM9URwCAx6we5ggpoLr/8u2Pms55
U0BQKKSIDG/hS3lb/XfPh+LP4rsB1FmJxCGsP8gmcizKIDspQw7kWVnxM70+Q/WL
1Ok5yQII7d0dd3IdOCGwARzlprsCepOTw5OiHMQFO8NwmeirV7vJzXWTU9eFAXIF
y7q4ZCw/Gxgy8f62/ag47y3HqUjJc2utpNTAnbLH2vqr1WZNFYK+WO3OM0br6xLV
JnRBdQuesHzJcXBal51u1LLeLpBcPtdNB613DMj7rYtxopjr8yTQgxmolrgE4YqU
vqpSrTFb1jlVN/IdgAVrGaCX53TfBSujMuyDpEO+HjOUd/KtAWK17c7ZbhVPtiiU
+wvIMkEAzROkybgKNc0gfA3Kxsnq24mgNXy53gjG3omdN5uXmfMsivl7iRI1yMdA
7VjojmdPiZS9z5AYrDrYXzx8g8FCE21OhD81CtRwagwRKXm/Pskc4yjbvMbjAMn/
34K484aUJgOE6pVRj9FwXRb7deN8uIRvOGWPueHxsg3i09yw8EOpnUboTxxgJ3hu
k/X/HXUTBGgVRmsce+iEMXKoH89vnlJBHeF+4NRVFleFqOck8NUxKDVuIYCTNkTN
W6fgib+8JFMdOnnLpPklPx5LUXhEQmNT5qrO9bHIN3Ejn4VNgL74CIVrNpmMl1DQ
`pragma protect end_protected
