// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:37 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fh54ibFfy/DzMr8gWRvzWi7CprJbrXKBdMjIcLEg0KKq0pd3OykoRscc+6rpOJTr
W105pyzBIvOEP4dqoZwdTsigP0kduWcdoNKlDl03o4GIH/rnTBP3XbeGs/hwd4FO
/JATVe9O/jT3y/wo93Mwayg0CPBNFzkkYlpLqP2uzUQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
eSVv74RFhwiVjsqvuy9JUVCb9XvW69D8Ql67kh5hEBN41VW1EcFVQ/QgIlC1pgue
hquW6WWCdTecOb1NHumAtiNlX9GxNoqC+t6IFMEXdPx7qpZDHkN4Reb9ZD0GyB3v
jWGOje/b4oUhRZ/6dhtk6s1PaCZDhKIMxq7bTfMcHeK/Xq86sOHiL8+gdOYZUGM3
77JmwAX7tju60AUMBz2jeMKh0rmSt7togoYdVO/MtqpMxWwuJ5gD4rUyacx5lWTO
2hP4v+jTO8gleTdMiGCjUGqZEBJONKpgziZCHifuDRN+MPl0xgwVZJeacv0Zwg+g
YHUba9fhFYPU5XVoln4iv7mquWM4MSnwO497GkRg1xEVOvbXu9rDqlmJMsIGqldJ
ZNEHmKJ7XtDxg/6d0Ni5TZ+RCx7JZHeEUavx4HqBuojaav3FYIuzS45UgK84iyJD
M3yMH30/BqPomN787Q1qUell74Lez6AcYUOPfRyR3bcF7tFhN02K1R2agvK5mIBA
ZaA4CKRWepIyWaiFPifEOwhYQILXhfPYUaMcRS5Splo9BIBDho9lcOi3OX7k4Wd4
HQXq2NFvslCAMuzEaYETg3eJiBw5RmikAEnF5YPIKFQb1QJ4Giz4vvpIPKoNvKdh
MEqihnMU8DMBX+XkPnNKVd+lM60m7GvX7nSmJg1LImvprv39l7e7vQK3xx2mbNkk
3w5/4sPjYYQ5ddzUVvxJqapXpdrqt7hBxzVzPTaEfv3xFa7jfn+1yTMJ/cgOImUk
dm1/3T6YSxOWBcQHSXK2eKdkZYSmdh6gx9/hBLI3yohO+0mTE3hBJUmDqnpxW2UM
fB8YD+1AbTJeg9SB5zeiQKOc+uIBhAkvdgmz501BPpYk5p0pw3tZLp3onLN2PknH
3ZSd+RpYbCaVA6JZGNz0aPRsAQFufVtV+8w8m0YEmpbAvq2DdTmJlNIi2y32nM39
d6+hZvlRTIq2UBROAYMFN8XY6bO8LgF4ZGa0zOglatjQi3zCtyMLXew5d+Jk/Fug
u8a2oF3dUFduaum1HPBUGAWc5nwaAgjBTK8SePiaWaanG+e6uuOUd6i5fV9aoywb
Qig1VFo3Kvt3W0mDjxIFYKCshdTLdPT/n9tWGuvQYo435jfcrluAQD+0XT5dM1Yu
C466+DyEw5DoAXHCVGq0OxZe8dYdp2oxc8UrdjfpCDVpY2INdmyORoiXvYKQuGN9
G76qFldJ8QYX2fNtDim+BWQcAycrInjRDdkDRMVL7Jl4DypNg86I1E+x7hof98/S
D2ammwdQAGrcdOrvGlhDp0xqG5ajmnLDEEX75veYZSbRtn2QQ0mE/wj5297UFTlB
263uJklUlniMsDLVRjj0726SCngfe7fu6oXaQiTH6xBzjm07PwdS5TakOCsDuhpR
XBIIJh8zKvIEl1qj15+XETlsJqwCOlfOhwQH0YCifU6avwujMvtpKHB3bQfjbsd+
Pc0pNsPZkZJLDGorBHXElOjfiEHKPMwkasC5Yj2h9YMwfLrumIsbF0tpIz5RSSGc
oHcNkfFbhRRpjkAMqXJ06lFogrph/loJ1HQuptdb++j1FOJ+z50Rtm9Hv0J/Lvke
ivBNwdRjJPMaJMm1L2ByGl+2svnNNkKm26z6XIBF7pP4WsDnJjQVtN6Eq6o6kuuO
Qc2xdfoYf8pbMqB9MOw6Hf2L7223/7nSFvvbHX4BWniaH/rZlmTPhS9hFFZFje5k
oGX8eGxJjX6FRm5daDELtIPGLcLBGmJsD6ayGbFUE2/Wuf9zMv690kZBy1QTO2Kh
3l5uN/VxAj8JMtVSJ0/OqvfyrN4YcaOOdluFcvqGhQu9+Lsm4TKTpW7vm+38kqnu
k3RpINXTf45EqG+GT5XPP6fmh0i/9c0PZ8JYEBW59Ud9sYr5ELizzCEgMeXeUeyg
Jw+x7SBdsVSrSJ1+8vJtgtaq1f1dqw7TetcbfICBh4kGgH/KvSCtVSmGdbI9vfM+
rP6MLYZdmN+GSk55AmPz050ZPt8gUhv2F8vJQObEbyHYwNsNbFQ9Qy3zY8rT2Y9f
OsjOMJnW400XgZAE7cwBhrZZ5dZpmCj/xAp1rOT6JG8k2m0Yp7vRSK0We4HqHIcu
XV8H+OhHftgkgOdWzAYOOisXgP71WyekiCDcs28XuRdILuh7P+5FWScG+mL25u8p
6ftPf1xGivy1L0YcWIpqvdH3HLt8HlzmEkEYSKkeutI7cSb2P3PGc++UCpzAG8wE
sLSTm/uuEcPoRa6lqixGkpmlPA2tJNxlelYN600Pq6h5dwnTATpfZygx2l8b7kWb
+uMkOSlV7YYJ/1w1d2lxAGgaP3UWqYZZLEPjw8VPWJirUZ6jpHXXZS36BdSiuB1a
XUlXODo0TOO1HV0lJhwbWSvA1OnyrwAJHUsvgF8uVRvVZkTPY7K/TabT7v5LPotI
jgSePPUXC3y5cKUVmFQwFqGSe0Yfet4xZjSn0Sw8xaE+EUaOAdMzAyUCRo9BRgqn
ZgMFzwZF+SFZ/TwRBhc4miSn3keZOICSle+Rk5RTtDVQtdJ+wL8LtGyPQNTYRPg1
B6uDt54OdnOusei+BKag6NDx+0/fiDJ3gjmwaiWcIAZ+LG5zM63DFQNh6oZ4Qdod
n1nkTZRY2Vn7xPhPqi5TpeNFWO6htZzmDnXKy4UcQFqO+j7vQcppN9dleAoom29j
jzHni9BRqVS2x5jygAgFlxKzT+bIFRIwBcxqrbpJbT/e1EOQLsbQSgHnEVqhUKDo
lHfn4q4tQieD7zo356Ms4tYM8fitxE9MIfzQ2ZC/CbTcO3yJ6DYYlojF7DXnH2le
VnliLyH2Bs2HHLcOPvYm3uXePA22KTicJBZgkmNl1TcRQ2FhNVJKZ9UyvD3OXS66
2VOfvEVyMwpFZEvTHYSzmSUuI3fMedSUxbJGl582bn61O9XT3yUc9n3sWpQutUXf
cv4uQKP365Ku/ajw5PXns4SUQ93qt/MKLAyp+j+rOOBhv1C9xF7SHCHIcGA6yGTV
ufpFNJl2mg8247dOMYUhX9SGCOE5hHBn70vySFKnHAKbJ3zpUo9zGCUyd2KldjMl
EY/tPjgkyt2d9eBqKdu5YmUGeWe7g51G3WiiIMKHs24CD2ktwvV2WWYQlyd4gRmX
/C32mS5JsH/Alb0D8gKq8DZyFTu9PVKgbq5bGSn0IGV+NEtmyphyTM7glYaZNU4a
+/A0ywv5ei15WM7WHJiNufjYAppSAqhjuLpJDApoAeF7Z/ixDCj8slS2ovcStu8c
veEqkc/ItqMXHWRpGF/5nzOaHWkKMiZUgIq8q+rz67ILnnkU4h51v8tycJ4b1ibx
2sKDzoCVoN3U4B6D9nesIqzSCSsE2kRyP4DqkQWcst785muBKUJqIAA3ELWanb74
D2uDYfmyHnrIrDJz3POY9ZAg6MnXk6GBnjloSG0vEqiG7s89f7xQjoGzYv/nccSe
Nq2653kn1gw4+lkdbWUmvVaGea50HQfM02QPEn971Qr//PTR7GKjELRI8PErl0go
Swson08Ga+UQ9cymMptnc+mR1xSqlmFJNH6xS0G5YUugUm/1pmcmRlnavyxuIYPv
3q3amw5IRnHXQ4Eoo1tMvqWB7+3wIFjkwqwAprzLp/WUcjslsr1h13H0x2K5pomF
VHoiCqD6fCp4NadkRvCEIZ3Blj3jbn19H5d4jms+fpvew78bOJh2Q2h/w8F+SE3b
LH5LsSssgKA0The+sdWYSG7hCyoFKtJhDW1xtbPO1rDuiJn9gffunyv/BJVcOooZ
qLiiLOyjuIu7vYqf36bhi0zgx3t7lFh8PA6SDAePk0BZeZcrJXbyz+pBfElKYUqk
jcJeeQHlHwSGwDB7Ii8ibhzjCDjhV0ZF8gEx5SlIQUCACyckLgX3bPSPQnhV3Rpa
tBsXsv3/ARK1NNUBofjW1nCa8fTqoe3IG1CYkYLg72ERA0FDJ4feOahcNEEeToLE
a4StVzZ96vgUNwlbXkfMCUnWDlmDBhwU7EA3VjbmoiTTjeTgsMBPBSv9M+Buxbah
sif5uGNnj2I7yvP+8ctZQCncaeFEtsD1UgK6Wj0SCLHN7Mz/MN8U/vgPN4wNvu3A
u79WcQZDT+2DNYKp3cT7COsruYkWC4fxqrEsBnamWW8oPqu5bCJ5dqxtPGg0f9Xg
rUVs6VbK4m18OALeSfDyfrXNhXvHA6jIC2q9NnT3Gi6dDI9jn+kJbkyfT1k4uvZX
Yx+eD4TgXo7TIhlx6Ng7luvaTvLCG76wJa8ju5HX3ofNnEB86lUmRIUNhAf7KaKq
pmmXeeITVTnkeVyPSPIIzQndp4RX6C+md32Odap2xoDsj6gSLKXNhqb4Hd2eQGt9
zVvX+GsotQi5FJfD63rm9ONCoLsTL8qvc7xGls0Hn2PbXHSkKeywxTO6zMj5wUpJ
E+WDeBkhA6qzEAIzErN4r8qEenTb9MGZUk8RmKcN92ejbCo+AbjKxYV7Io/4z6bp
wr7SrxX1PSTFw7nZ6l7pxhNa+BFvMW/SaX0EPX204WbLZ589n7p11aYcm1kSKKe5
VAtASfbBPdlmlC/sfU9D0L7uFBSVOgdg9jjKU9oeNmLVzhmB8ejBIXLeEY/e3Rds
c3GXhGJqTIDFsjJfz3ujEoEkMY0cM0QuGSzxU4hjSPsxtGWd6TjRO1xTopLtdrjQ
Z3jRYZh73WIT4gWEa/7azwlqaikwcqwSyq/4zzhS7my+gp75+klMxbc9kXUJpeP+
GGGMetO0cTInuCxgto8QNJyD78uez4dAvKZgp41iu3m0utNOdk7oQ+bGvVk/CZfi
Iup3PIxcc3x8wYkCGDNDsyxtug5GyfJlZIJjxYPqVgxdbn5keILFU30sFv0IiFkR
9R7VlbPeossG6SABXuSsKOQMbriMQgtwcSOq/xXKLa49XsKWvPVLToELyNFPPgem
7G23N7XAGkqoezzwGWWJ/em6B9GP3vKPgBINJaeywTFJcJgsB2+pde4qPJNdB7iS
k8vNC0wLRaAsTp5GTuJ7x4VNQ4Hp4DLHNmL680rlvBS9q57wOvkUVY+7dSd6omk3
Lycos8Kq9l1N9CMVAu4J7MZO+EPwJi/BPkcuj757kCTNd56qjvhxyJFPWrIK5tx7
FwD5nNMtyhe/UfwFD9Yeo0EdkneDccz/ZQlzNsoZfjgbO6ewWJ5nkdanY/mPxXNT
elrus3lJnCH+nBtpSNb9OU75kAvyNrYCXdo+n03unaOUBvp+Z121V7Hx3gorXfVU
aB32iXVMEKl0Q51N9RHRWFp/UonPCiZ4tVOViZ+ZrlPxQWGbEL2RLCgOCQOCI4bL
fE/fQQTlSpIZwVCDNmh5UUNBAmXJJft8IjErmzz3Z3XA6WaCQj8xKkjSI/eRxdhM
bNB9YvUjSkrAfGZMMBGcRS7ZI4eG6i+D9YXqQIxccP/mVyNBRQWp622ST0TSFE4f
11dI9kT/54ByEAxgYsD7uqd9/NEkinGinVFNhdC0zkuxrHlV/aFx4kYYH3amPvIY
5Zg1a0xPwqHwoihftzjfIKT71OxtH8EN+xJsLcDQD2nXC28mLJGrUgrDyrEz0W6X
XyBvOJdm9XRTZkCsyiJYU2l/3USYfNDZ2KT3lL22b94KEFINamCfvGmukKCd8SSG
gGLhY2KFvrKzMeGAlFaOUKKYRLQmzD6INs7sLeObmxxvf7KCfUJoxYM5XP0+hAPX
p4yfqlO4h2Ln4IdYm/LnN1Zsfi9b1DpIqPvd4evEeEbBla7wv7elPP6/+35sKAhU
fhRvxvwFzZ1shlqYpWdCQE5F3RQ7z7I8wceRDegPXnZg023oSNhZmaqbRHd/AltL
ku6SzLJw76xSNxSfhGJEjfO+KjDkYFz9m9syXAq2eI5hkVPthkDk/r8ywA8UpmlK
XlHPFlgFhx4E08rRbyUehkCxrK1aAygWG8UjjClbBlqnWT48AuMPN8EPX6MSe8na
X5xdR2xAiNHiHYY2j9GsSTwasn1hVw2BAP71sXuJT6WmA0vAyKjZEok/b+rg0zwg
jn0QhPUOp7AlUKr4jqEeliW8vndQS2XNl6ASCXKHt0ztQ/H65YVtENZEA7LdT0Kp
gJ5E/iHPJyLcZCTDhWtF9SM9fXzF5bAUXBAkg2n65Xu0XBbAwDbdZBbGeAvgzZ+k
e7+TxInl1FRDGXfYYf8KDqNmGfyi4DtRI273Sepy0cjHllE/0xZryNR7xK9JlztI
YxLNWQE9JU1vbxRp3dFjoKX5jDU0eYR568yua8qFhE9kZSvtg2VPRwHY8ES0bEFG
5LdB55F7q7LeMo77eARbGV12WdjrJvKqtJf6vfi7Mj7HphU7Wn0K38Jn7lHYxnLG
iTLF/h9ZzT2OdnoZweNvnttKe3InOmIg7gc6xzSYizu2zTv9jJSYdRKv9v8NtCAd
jWIPCD1mlQmjIunFaaE41qBTUIGHPdlcF4hA5z0q3pCm7AeFFhoW9c12oZH7XfrG
cqMSCcp37dSNdQYF3A5Flw+eL1tP+VrAJt50kFpqQU5u7P8CM2jW57G89dkJF4JY
QeRUwCxYisSjFL/olDt8DlfqFxAzjI9rJWItUAZZ+6fKMNRmhvMYqnR9SSO19y+/
o+HjvGAeYUbzx5SGwNZRtOTggWWgJMJif3PaSD+brekDOz4w11ZcBYUbeIomItLM
Vs+WmP+jqfIq18XtPFvO/RmXVdk5LFkXEdfC5inQvil3X5wTYz3UjXOswoyrvrL2
bnC90yBjl5JULtzsHw9b12P/9OiZ4J8NG48u3LlcFgCi+ony3kQPB1BJ/YziYfte
gEoevHTj5LFUxEJxU6n9AkRJ/wH62cOdhNYMGL7AFP3fy0XOT/Oiw6YXKFOAbuEW
UB/ksZCbQCO5C9pAPJA7AMD1Aw7GF/bW42vhuq8hbs6dL8oDLbNvuyjnXgHkugTd
HKut/2yR/JT27WZ1BNBG+0/vsrY6V6IcRfn5KNRyffctKyEbpk1r+BdY6H4DwMUT
NWxdqa0q1UeZv9KLFwQrXrTGSQEeB8zN0poouCjcQloe0/tCilQwf/8Zbno5CQpo
kxEnFiIiTMbOtKMSMqUgexF94kv0aPQM38eprMV08Yqq42DFNc5pIyH7qflFpdwE
SuChqesvQAr+a6qRdR2CV3EFA3xHc9mZzi7BPnT8OGR0Y3D7R8CNSd5VqmrruxPP
s0KOjmBoJRoU5QBmLl+AWxg+WVuaqzawUnf7Yq8uXGyBh6f6sv1cuwvZHOFaiZVO
qngHcKrLUypevI45kx4RVWlnkUqCp52JjUmkbf04NvCExAqZRtG3HXaX/sH+EApd
OSF+FLURXL7nssJgvltZ6bl44xr5pJV9iLYzFzmquu9I1kQbQTJx1WDh2zZI5htT
oGaPsNc96Vr0f1oGj9rDtKgCxB3X+qqG/Jn9hP7nYzveOuM1eoEcB8wn5p74cj5F
GKNv9KqEToOxyChcqWO5/tpiMKQ/qaFjtOZrdqLt+KcN0ScLQw7ffpZCYvoGK2Gk
qev25pOTJN17hh84nTeUvTBJnExZvLVzjf1TgVTA7eH2QuMZM2VEH5IuFP8VblYK
q9v9RUr0yStV7UJcT7yY58bV+adkJTxUgYIOfhpw7toOt/v6prs+8+sW8+4tsAHe
w7yLGJC2n203H3tS5ERrIQ==
`pragma protect end_protected
