// pcie_cv_qsys.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module pcie_cv_qsys (
		input  wire        clk_clk,                                                //                                    clk.clk
		input  wire [31:0] pcie_cv_hip_avmm_0_hip_ctrl_test_in,                    //            pcie_cv_hip_avmm_0_hip_ctrl.test_in
		input  wire        pcie_cv_hip_avmm_0_hip_ctrl_simu_mode_pipe,             //                                       .simu_mode_pipe
		input  wire        pcie_cv_hip_avmm_0_hip_serial_rx_in0,                   //          pcie_cv_hip_avmm_0_hip_serial.rx_in0
		input  wire        pcie_cv_hip_avmm_0_hip_serial_rx_in1,                   //                                       .rx_in1
		input  wire        pcie_cv_hip_avmm_0_hip_serial_rx_in2,                   //                                       .rx_in2
		input  wire        pcie_cv_hip_avmm_0_hip_serial_rx_in3,                   //                                       .rx_in3
		output wire        pcie_cv_hip_avmm_0_hip_serial_tx_out0,                  //                                       .tx_out0
		output wire        pcie_cv_hip_avmm_0_hip_serial_tx_out1,                  //                                       .tx_out1
		output wire        pcie_cv_hip_avmm_0_hip_serial_tx_out2,                  //                                       .tx_out2
		output wire        pcie_cv_hip_avmm_0_hip_serial_tx_out3,                  //                                       .tx_out3
		input  wire        pcie_cv_hip_avmm_0_npor_npor,                           //                pcie_cv_hip_avmm_0_npor.npor
		input  wire        pcie_cv_hip_avmm_0_npor_pin_perst,                      //                                       .pin_perst
		output wire        pcie_cv_hip_avmm_0_nreset_status_reset_n,               //       pcie_cv_hip_avmm_0_nreset_status.reset_n
		output wire        pcie_cv_hip_avmm_0_reconfig_clk_locked_fixedclk_locked, // pcie_cv_hip_avmm_0_reconfig_clk_locked.fixedclk_locked
		input  wire        reset_reset_n                                           //                                  reset.reset_n
	);

	wire          pcie_cv_hip_avmm_0_coreclkout_clk;                               // pcie_cv_hip_avmm_0:coreclkout -> [irq_mapper:clk, mm_interconnect_0:pcie_cv_hip_avmm_0_coreclkout_clk, mm_interconnect_1:pcie_cv_hip_avmm_0_coreclkout_clk, mm_interconnect_2:pcie_cv_hip_avmm_0_coreclkout_clk, onchip_memory2_0:clk, rst_controller_001:clk, rst_controller_002:clk]
	wire          alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy;                 // alt_xcvr_reconfig_0:reconfig_busy -> pcie_cv_hip_avmm_0:busy_xcvr_reconfig
	wire  [229:0] pcie_cv_hip_avmm_0_reconfig_from_xcvr_reconfig_from_xcvr;        // pcie_cv_hip_avmm_0:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [349:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr;           // alt_xcvr_reconfig_0:reconfig_to_xcvr -> pcie_cv_hip_avmm_0:reconfig_to_xcvr
	wire          pcie_cv_hip_avmm_0_rxm_bar0_waitrequest;                         // mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_waitrequest -> pcie_cv_hip_avmm_0:RxmWaitRequest_0_i
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar0_readdata;                            // mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_readdata -> pcie_cv_hip_avmm_0:RxmReadData_0_i
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar0_address;                             // pcie_cv_hip_avmm_0:RxmAddress_0_o -> mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_address
	wire          pcie_cv_hip_avmm_0_rxm_bar0_read;                                // pcie_cv_hip_avmm_0:RxmRead_0_o -> mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_read
	wire    [7:0] pcie_cv_hip_avmm_0_rxm_bar0_byteenable;                          // pcie_cv_hip_avmm_0:RxmByteEnable_0_o -> mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_byteenable
	wire          pcie_cv_hip_avmm_0_rxm_bar0_readdatavalid;                       // mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_readdatavalid -> pcie_cv_hip_avmm_0:RxmReadDataValid_0_i
	wire          pcie_cv_hip_avmm_0_rxm_bar0_write;                               // pcie_cv_hip_avmm_0:RxmWrite_0_o -> mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_write
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar0_writedata;                           // pcie_cv_hip_avmm_0:RxmWriteData_0_o -> mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_writedata
	wire    [6:0] pcie_cv_hip_avmm_0_rxm_bar0_burstcount;                          // pcie_cv_hip_avmm_0:RxmBurstCount_0_o -> mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_burstcount
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;                // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                  // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire    [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                   // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire    [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;                     // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                 // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;                     // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire          pcie_cv_hip_avmm_0_rxm_bar2_waitrequest;                         // mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_waitrequest -> pcie_cv_hip_avmm_0:RxmWaitRequest_2_i
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar2_readdata;                            // mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_readdata -> pcie_cv_hip_avmm_0:RxmReadData_2_i
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar2_address;                             // pcie_cv_hip_avmm_0:RxmAddress_2_o -> mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_address
	wire          pcie_cv_hip_avmm_0_rxm_bar2_read;                                // pcie_cv_hip_avmm_0:RxmRead_2_o -> mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_read
	wire    [7:0] pcie_cv_hip_avmm_0_rxm_bar2_byteenable;                          // pcie_cv_hip_avmm_0:RxmByteEnable_2_o -> mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_byteenable
	wire          pcie_cv_hip_avmm_0_rxm_bar2_readdatavalid;                       // mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_readdatavalid -> pcie_cv_hip_avmm_0:RxmReadDataValid_2_i
	wire          pcie_cv_hip_avmm_0_rxm_bar2_write;                               // pcie_cv_hip_avmm_0:RxmWrite_2_o -> mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_write
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar2_writedata;                           // pcie_cv_hip_avmm_0:RxmWriteData_2_o -> mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_writedata
	wire    [6:0] pcie_cv_hip_avmm_0_rxm_bar2_burstcount;                          // pcie_cv_hip_avmm_0:RxmBurstCount_2_o -> mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_burstcount
	wire   [31:0] mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_readdata;    // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> mm_interconnect_1:alt_xcvr_reconfig_0_reconfig_mgmt_readdata
	wire          mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest; // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> mm_interconnect_1:alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest
	wire    [6:0] mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_address;     // mm_interconnect_1:alt_xcvr_reconfig_0_reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_read;        // mm_interconnect_1:alt_xcvr_reconfig_0_reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire          mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_write;       // mm_interconnect_1:alt_xcvr_reconfig_0_reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire   [31:0] mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_writedata;   // mm_interconnect_1:alt_xcvr_reconfig_0_reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire          pcie_cv_hip_avmm_0_rxm_bar4_waitrequest;                         // mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_waitrequest -> pcie_cv_hip_avmm_0:RxmWaitRequest_4_i
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar4_readdata;                            // mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_readdata -> pcie_cv_hip_avmm_0:RxmReadData_4_i
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar4_address;                             // pcie_cv_hip_avmm_0:RxmAddress_4_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_address
	wire          pcie_cv_hip_avmm_0_rxm_bar4_read;                                // pcie_cv_hip_avmm_0:RxmRead_4_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_read
	wire    [7:0] pcie_cv_hip_avmm_0_rxm_bar4_byteenable;                          // pcie_cv_hip_avmm_0:RxmByteEnable_4_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_byteenable
	wire          pcie_cv_hip_avmm_0_rxm_bar4_readdatavalid;                       // mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_readdatavalid -> pcie_cv_hip_avmm_0:RxmReadDataValid_4_i
	wire          pcie_cv_hip_avmm_0_rxm_bar4_write;                               // pcie_cv_hip_avmm_0:RxmWrite_4_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_write
	wire   [63:0] pcie_cv_hip_avmm_0_rxm_bar4_writedata;                           // pcie_cv_hip_avmm_0:RxmWriteData_4_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_writedata
	wire    [6:0] pcie_cv_hip_avmm_0_rxm_bar4_burstcount;                          // pcie_cv_hip_avmm_0:RxmBurstCount_4_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_burstcount
	wire          mm_interconnect_2_pcie_cv_hip_avmm_0_cra_chipselect;             // mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_chipselect -> pcie_cv_hip_avmm_0:CraChipSelect_i
	wire   [31:0] mm_interconnect_2_pcie_cv_hip_avmm_0_cra_readdata;               // pcie_cv_hip_avmm_0:CraReadData_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_readdata
	wire          mm_interconnect_2_pcie_cv_hip_avmm_0_cra_waitrequest;            // pcie_cv_hip_avmm_0:CraWaitRequest_o -> mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_waitrequest
	wire   [13:0] mm_interconnect_2_pcie_cv_hip_avmm_0_cra_address;                // mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_address -> pcie_cv_hip_avmm_0:CraAddress_i
	wire          mm_interconnect_2_pcie_cv_hip_avmm_0_cra_read;                   // mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_read -> pcie_cv_hip_avmm_0:CraRead
	wire    [3:0] mm_interconnect_2_pcie_cv_hip_avmm_0_cra_byteenable;             // mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_byteenable -> pcie_cv_hip_avmm_0:CraByteEnable_i
	wire          mm_interconnect_2_pcie_cv_hip_avmm_0_cra_write;                  // mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_write -> pcie_cv_hip_avmm_0:CraWrite
	wire   [31:0] mm_interconnect_2_pcie_cv_hip_avmm_0_cra_writedata;              // mm_interconnect_2:pcie_cv_hip_avmm_0_Cra_writedata -> pcie_cv_hip_avmm_0:CraWriteData_i
	wire          irq_mapper_receiver0_irq;                                        // pcie_cv_hip_avmm_0:CraIrq_o -> irq_mapper:receiver0_irq
	wire   [15:0] pcie_cv_hip_avmm_0_rxmirq_irq;                                   // irq_mapper:sender_irq -> pcie_cv_hip_avmm_0:RxmIrq_i
	wire          rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, mm_interconnect_1:alt_xcvr_reconfig_0_mgmt_rst_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	wire          rst_controller_001_reset_out_reset_req;                          // rst_controller_001:reset_req -> onchip_memory2_0:reset_req
	wire          rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:pcie_cv_hip_avmm_0_Rxm_BAR0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pcie_cv_hip_avmm_0_Rxm_BAR2_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:pcie_cv_hip_avmm_0_Rxm_BAR4_translator_reset_reset_bridge_in_reset_reset]

	alt_xcvr_reconfig #(
		.device_family                 ("Cyclone V"),
		.number_of_reconfig_interfaces (5),
		.enable_offset                 (1),
		.enable_lc                     (0),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (0),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),                 //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_clk),                                                         //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                                  //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_address),     //      reconfig_mgmt.address
		.reconfig_mgmt_read        (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_read),        //                   .read
		.reconfig_mgmt_readdata    (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_readdata),    //                   .readdata
		.reconfig_mgmt_waitrequest (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest), //                   .waitrequest
		.reconfig_mgmt_write       (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_write),       //                   .write
		.reconfig_mgmt_writedata   (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_writedata),   //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),           //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie_cv_hip_avmm_0_reconfig_from_xcvr_reconfig_from_xcvr),        // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                                //        (terminated)
		.rx_cal_busy               (),                                                                //        (terminated)
		.cal_busy_in               (1'b0),                                                            //        (terminated)
		.reconfig_mif_address      (),                                                                //        (terminated)
		.reconfig_mif_read         (),                                                                //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                            //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                             //        (terminated)
	);

	pcie_cv_qsys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pcie_cv_hip_avmm_0_coreclkout_clk),                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	altpcie_cv_hip_avmm_hwtcl #(
		.lane_mask_hwtcl                          ("x4"),
		.gen123_lane_rate_mode_hwtcl              ("Gen1 (2.5 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.in_cvp_mode_hwtcl                        (0),
		.bar0_size_mask_hwtcl                     (12),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Enabled"),
		.bar0_prefetchable_hwtcl                  ("Enabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (9),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Enabled"),
		.bar2_prefetchable_hwtcl                  ("Enabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (14),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Enabled"),
		.bar4_prefetchable_hwtcl                  ("Enabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.CB_P2A_AVALON_ADDR_B0                    (0),
		.CB_P2A_AVALON_ADDR_B1                    (0),
		.CB_P2A_AVALON_ADDR_B2                    (0),
		.CB_P2A_AVALON_ADDR_B3                    (0),
		.CB_P2A_AVALON_ADDR_B4                    (0),
		.CB_P2A_AVALON_ADDR_B5                    (0),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (57353),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (0),
		.subsystem_vendor_id_hwtcl                (0),
		.subsystem_device_id_hwtcl                (0),
		.max_payload_size_hwtcl                   (128),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.rx_ei_l0s_hwtcl                          (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (4466),
		.vsec_rev_hwtcl                           (0),
		.user_id_hwtcl                            (0),
		.avmm_width_hwtcl                         (64),
		.AVALON_ADDR_WIDTH                        (64),
		.avmm_burst_width_hwtcl                   (7),
		.CB_PCIE_MODE                             (0),
		.CB_PCIE_RX_LITE                          (0),
		.CB_RXM_DATA_WIDTH                        (64),
		.CG_AVALON_S_ADDR_WIDTH                   (32),
		.CG_IMPL_CRA_AV_SLAVE_PORT                (1),
		.CG_ENABLE_ADVANCED_INTERRUPT             (0),
		.CG_ENABLE_A2P_INTERRUPT                  (0),
		.CB_A2P_ADDR_MAP_IS_FIXED                 (0),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES              (2),
		.BYPASSS_A2P_TRANSLATION                  (0),
		.a2p_pass_thru_bits                       (8),
		.ast_width_hwtcl                          ("Avalon-ST 64-bit"),
		.use_ast_parity                           (0),
		.reconfig_to_xcvr_width                   (350),
		.hip_hard_reset_hwtcl                     (1),
		.reconfig_from_xcvr_width                 (230),
		.bypass_cdc_hwtcl                         ("false"),
		.single_rx_detect_hwtcl                   (4),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.maximum_current_hwtcl                    (0),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l0s_aspm_hwtcl                    ("true"),
		.extended_tag_reset_hwtcl                 ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.aspm_config_management_hwtcl             ("false"),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("true"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     (0),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.millisecond_cycle_count_hwtcl            (124250),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (67),
		.cpl_spc_data_hwtcl                       (269),
		.coreclkout_hip_phaseshift_hwtcl          ("0 ps"),
		.pldclk_hip_phase_shift_hwtcl             ("0 ps"),
		.port_width_be_hwtcl                      (8),
		.port_width_data_hwtcl                    (64),
		.hip_reconfig_hwtcl                       (0),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_clk_switch_hwtcl                  ("disable"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.no_command_completed_hwtcl               ("false"),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.deemphasis_enable_hwtcl                  ("false"),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("true"),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (255),
		.reserved_debug_hwtcl                     (0),
		.use_tl_cfg_sync_hwtcl                    (1),
		.diffclock_nfts_count_hwtcl               (255),
		.sameclock_nfts_count_hwtcl               (255),
		.l2_async_logic_hwtcl                     ("disable"),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.indicator_hwtcl                          (0),
		.rpre_emph_a_val_hwtcl                    (11),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (22),
		.rpre_emph_d_val_hwtcl                    (12),
		.rpre_emph_e_val_hwtcl                    (21),
		.rvod_sel_a_val_hwtcl                     (50),
		.rvod_sel_b_val_hwtcl                     (34),
		.rvod_sel_c_val_hwtcl                     (50),
		.rvod_sel_d_val_hwtcl                     (50),
		.rvod_sel_e_val_hwtcl                     (9)
	) pcie_cv_hip_avmm_0 (
		.coreclkout           (pcie_cv_hip_avmm_0_coreclkout_clk),                        //          coreclkout.clk
		.refclk               (clk_clk),                                                  //              refclk.clk
		.npor                 (pcie_cv_hip_avmm_0_npor_npor),                             //                npor.npor
		.pin_perst            (pcie_cv_hip_avmm_0_npor_pin_perst),                        //                    .pin_perst
		.reset_status         (pcie_cv_hip_avmm_0_nreset_status_reset_n),                 //       nreset_status.reset_n
		.test_in              (pcie_cv_hip_avmm_0_hip_ctrl_test_in),                      //            hip_ctrl.test_in
		.simu_mode_pipe       (pcie_cv_hip_avmm_0_hip_ctrl_simu_mode_pipe),               //                    .simu_mode_pipe
		.RxmAddress_0_o       (pcie_cv_hip_avmm_0_rxm_bar0_address),                      //            Rxm_BAR0.address
		.RxmRead_0_o          (pcie_cv_hip_avmm_0_rxm_bar0_read),                         //                    .read
		.RxmWaitRequest_0_i   (pcie_cv_hip_avmm_0_rxm_bar0_waitrequest),                  //                    .waitrequest
		.RxmWrite_0_o         (pcie_cv_hip_avmm_0_rxm_bar0_write),                        //                    .write
		.RxmReadDataValid_0_i (pcie_cv_hip_avmm_0_rxm_bar0_readdatavalid),                //                    .readdatavalid
		.RxmReadData_0_i      (pcie_cv_hip_avmm_0_rxm_bar0_readdata),                     //                    .readdata
		.RxmWriteData_0_o     (pcie_cv_hip_avmm_0_rxm_bar0_writedata),                    //                    .writedata
		.RxmBurstCount_0_o    (pcie_cv_hip_avmm_0_rxm_bar0_burstcount),                   //                    .burstcount
		.RxmByteEnable_0_o    (pcie_cv_hip_avmm_0_rxm_bar0_byteenable),                   //                    .byteenable
		.RxmAddress_2_o       (pcie_cv_hip_avmm_0_rxm_bar2_address),                      //            Rxm_BAR2.address
		.RxmRead_2_o          (pcie_cv_hip_avmm_0_rxm_bar2_read),                         //                    .read
		.RxmWaitRequest_2_i   (pcie_cv_hip_avmm_0_rxm_bar2_waitrequest),                  //                    .waitrequest
		.RxmWrite_2_o         (pcie_cv_hip_avmm_0_rxm_bar2_write),                        //                    .write
		.RxmReadDataValid_2_i (pcie_cv_hip_avmm_0_rxm_bar2_readdatavalid),                //                    .readdatavalid
		.RxmReadData_2_i      (pcie_cv_hip_avmm_0_rxm_bar2_readdata),                     //                    .readdata
		.RxmWriteData_2_o     (pcie_cv_hip_avmm_0_rxm_bar2_writedata),                    //                    .writedata
		.RxmBurstCount_2_o    (pcie_cv_hip_avmm_0_rxm_bar2_burstcount),                   //                    .burstcount
		.RxmByteEnable_2_o    (pcie_cv_hip_avmm_0_rxm_bar2_byteenable),                   //                    .byteenable
		.RxmAddress_4_o       (pcie_cv_hip_avmm_0_rxm_bar4_address),                      //            Rxm_BAR4.address
		.RxmRead_4_o          (pcie_cv_hip_avmm_0_rxm_bar4_read),                         //                    .read
		.RxmWaitRequest_4_i   (pcie_cv_hip_avmm_0_rxm_bar4_waitrequest),                  //                    .waitrequest
		.RxmWrite_4_o         (pcie_cv_hip_avmm_0_rxm_bar4_write),                        //                    .write
		.RxmReadDataValid_4_i (pcie_cv_hip_avmm_0_rxm_bar4_readdatavalid),                //                    .readdatavalid
		.RxmReadData_4_i      (pcie_cv_hip_avmm_0_rxm_bar4_readdata),                     //                    .readdata
		.RxmWriteData_4_o     (pcie_cv_hip_avmm_0_rxm_bar4_writedata),                    //                    .writedata
		.RxmBurstCount_4_o    (pcie_cv_hip_avmm_0_rxm_bar4_burstcount),                   //                    .burstcount
		.RxmByteEnable_4_o    (pcie_cv_hip_avmm_0_rxm_bar4_byteenable),                   //                    .byteenable
		.RxmIrq_i             (pcie_cv_hip_avmm_0_rxmirq_irq),                            //              RxmIrq.irq
		.reconfig_to_xcvr     (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),    //    reconfig_to_xcvr.reconfig_to_xcvr
		.busy_xcvr_reconfig   (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),          //       reconfig_busy.reconfig_busy
		.reconfig_from_xcvr   (pcie_cv_hip_avmm_0_reconfig_from_xcvr_reconfig_from_xcvr), //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (pcie_cv_hip_avmm_0_reconfig_clk_locked_fixedclk_locked),   // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (pcie_cv_hip_avmm_0_hip_serial_rx_in0),                     //          hip_serial.rx_in0
		.rx_in1               (pcie_cv_hip_avmm_0_hip_serial_rx_in1),                     //                    .rx_in1
		.rx_in2               (pcie_cv_hip_avmm_0_hip_serial_rx_in2),                     //                    .rx_in2
		.rx_in3               (pcie_cv_hip_avmm_0_hip_serial_rx_in3),                     //                    .rx_in3
		.tx_out0              (pcie_cv_hip_avmm_0_hip_serial_tx_out0),                    //                    .tx_out0
		.tx_out1              (pcie_cv_hip_avmm_0_hip_serial_tx_out1),                    //                    .tx_out1
		.tx_out2              (pcie_cv_hip_avmm_0_hip_serial_tx_out2),                    //                    .tx_out2
		.tx_out3              (pcie_cv_hip_avmm_0_hip_serial_tx_out3),                    //                    .tx_out3
		.sim_pipe_pclk_in     (),                                                         //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (),                                                         //                    .sim_pipe_rate
		.sim_ltssmstate       (),                                                         //                    .sim_ltssmstate
		.eidleinfersel0       (),                                                         //                    .eidleinfersel0
		.eidleinfersel1       (),                                                         //                    .eidleinfersel1
		.eidleinfersel2       (),                                                         //                    .eidleinfersel2
		.eidleinfersel3       (),                                                         //                    .eidleinfersel3
		.powerdown0           (),                                                         //                    .powerdown0
		.powerdown1           (),                                                         //                    .powerdown1
		.powerdown2           (),                                                         //                    .powerdown2
		.powerdown3           (),                                                         //                    .powerdown3
		.rxpolarity0          (),                                                         //                    .rxpolarity0
		.rxpolarity1          (),                                                         //                    .rxpolarity1
		.rxpolarity2          (),                                                         //                    .rxpolarity2
		.rxpolarity3          (),                                                         //                    .rxpolarity3
		.txcompl0             (),                                                         //                    .txcompl0
		.txcompl1             (),                                                         //                    .txcompl1
		.txcompl2             (),                                                         //                    .txcompl2
		.txcompl3             (),                                                         //                    .txcompl3
		.txdata0              (),                                                         //                    .txdata0
		.txdata1              (),                                                         //                    .txdata1
		.txdata2              (),                                                         //                    .txdata2
		.txdata3              (),                                                         //                    .txdata3
		.txdatak0             (),                                                         //                    .txdatak0
		.txdatak1             (),                                                         //                    .txdatak1
		.txdatak2             (),                                                         //                    .txdatak2
		.txdatak3             (),                                                         //                    .txdatak3
		.txdetectrx0          (),                                                         //                    .txdetectrx0
		.txdetectrx1          (),                                                         //                    .txdetectrx1
		.txdetectrx2          (),                                                         //                    .txdetectrx2
		.txdetectrx3          (),                                                         //                    .txdetectrx3
		.txelecidle0          (),                                                         //                    .txelecidle0
		.txelecidle1          (),                                                         //                    .txelecidle1
		.txelecidle2          (),                                                         //                    .txelecidle2
		.txelecidle3          (),                                                         //                    .txelecidle3
		.txswing0             (),                                                         //                    .txswing0
		.txswing1             (),                                                         //                    .txswing1
		.txswing2             (),                                                         //                    .txswing2
		.txswing3             (),                                                         //                    .txswing3
		.txmargin0            (),                                                         //                    .txmargin0
		.txmargin1            (),                                                         //                    .txmargin1
		.txmargin2            (),                                                         //                    .txmargin2
		.txmargin3            (),                                                         //                    .txmargin3
		.txdeemph0            (),                                                         //                    .txdeemph0
		.txdeemph1            (),                                                         //                    .txdeemph1
		.txdeemph2            (),                                                         //                    .txdeemph2
		.txdeemph3            (),                                                         //                    .txdeemph3
		.phystatus0           (),                                                         //                    .phystatus0
		.phystatus1           (),                                                         //                    .phystatus1
		.phystatus2           (),                                                         //                    .phystatus2
		.phystatus3           (),                                                         //                    .phystatus3
		.rxdata0              (),                                                         //                    .rxdata0
		.rxdata1              (),                                                         //                    .rxdata1
		.rxdata2              (),                                                         //                    .rxdata2
		.rxdata3              (),                                                         //                    .rxdata3
		.rxdatak0             (),                                                         //                    .rxdatak0
		.rxdatak1             (),                                                         //                    .rxdatak1
		.rxdatak2             (),                                                         //                    .rxdatak2
		.rxdatak3             (),                                                         //                    .rxdatak3
		.rxelecidle0          (),                                                         //                    .rxelecidle0
		.rxelecidle1          (),                                                         //                    .rxelecidle1
		.rxelecidle2          (),                                                         //                    .rxelecidle2
		.rxelecidle3          (),                                                         //                    .rxelecidle3
		.rxstatus0            (),                                                         //                    .rxstatus0
		.rxstatus1            (),                                                         //                    .rxstatus1
		.rxstatus2            (),                                                         //                    .rxstatus2
		.rxstatus3            (),                                                         //                    .rxstatus3
		.rxvalid0             (),                                                         //                    .rxvalid0
		.rxvalid1             (),                                                         //                    .rxvalid1
		.rxvalid2             (),                                                         //                    .rxvalid2
		.rxvalid3             (),                                                         //                    .rxvalid3
		.TxsChipSelect_i      (),                                                         //                 Txs.chipselect
		.TxsByteEnable_i      (),                                                         //                    .byteenable
		.TxsReadData_o        (),                                                         //                    .readdata
		.TxsWriteData_i       (),                                                         //                    .writedata
		.TxsRead_i            (),                                                         //                    .read
		.TxsWrite_i           (),                                                         //                    .write
		.TxsBurstCount_i      (),                                                         //                    .burstcount
		.TxsReadDataValid_o   (),                                                         //                    .readdatavalid
		.TxsWaitRequest_o     (),                                                         //                    .waitrequest
		.TxsAddress_i         (),                                                         //                    .address
		.CraChipSelect_i      (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_chipselect),      //                 Cra.chipselect
		.CraAddress_i         (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_address),         //                    .address
		.CraByteEnable_i      (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_byteenable),      //                    .byteenable
		.CraRead              (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_read),            //                    .read
		.CraReadData_o        (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_readdata),        //                    .readdata
		.CraWrite             (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_write),           //                    .write
		.CraWriteData_i       (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_writedata),       //                    .writedata
		.CraWaitRequest_o     (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_waitrequest),     //                    .waitrequest
		.CraIrq_o             (irq_mapper_receiver0_irq),                                 //              CraIrq.irq
		.rx_in4               (1'b0),                                                     //         (terminated)
		.rx_in5               (1'b0),                                                     //         (terminated)
		.rx_in6               (1'b0),                                                     //         (terminated)
		.rx_in7               (1'b0),                                                     //         (terminated)
		.tx_out4              (),                                                         //         (terminated)
		.tx_out5              (),                                                         //         (terminated)
		.tx_out6              (),                                                         //         (terminated)
		.tx_out7              (),                                                         //         (terminated)
		.eidleinfersel4       (),                                                         //         (terminated)
		.eidleinfersel5       (),                                                         //         (terminated)
		.eidleinfersel6       (),                                                         //         (terminated)
		.eidleinfersel7       (),                                                         //         (terminated)
		.powerdown4           (),                                                         //         (terminated)
		.powerdown5           (),                                                         //         (terminated)
		.powerdown6           (),                                                         //         (terminated)
		.powerdown7           (),                                                         //         (terminated)
		.rxpolarity4          (),                                                         //         (terminated)
		.rxpolarity5          (),                                                         //         (terminated)
		.rxpolarity6          (),                                                         //         (terminated)
		.rxpolarity7          (),                                                         //         (terminated)
		.txcompl4             (),                                                         //         (terminated)
		.txcompl5             (),                                                         //         (terminated)
		.txcompl6             (),                                                         //         (terminated)
		.txcompl7             (),                                                         //         (terminated)
		.txdata4              (),                                                         //         (terminated)
		.txdata5              (),                                                         //         (terminated)
		.txdata6              (),                                                         //         (terminated)
		.txdata7              (),                                                         //         (terminated)
		.txdatak4             (),                                                         //         (terminated)
		.txdatak5             (),                                                         //         (terminated)
		.txdatak6             (),                                                         //         (terminated)
		.txdatak7             (),                                                         //         (terminated)
		.txdetectrx4          (),                                                         //         (terminated)
		.txdetectrx5          (),                                                         //         (terminated)
		.txdetectrx6          (),                                                         //         (terminated)
		.txdetectrx7          (),                                                         //         (terminated)
		.txelecidle4          (),                                                         //         (terminated)
		.txelecidle5          (),                                                         //         (terminated)
		.txelecidle6          (),                                                         //         (terminated)
		.txelecidle7          (),                                                         //         (terminated)
		.txswing4             (),                                                         //         (terminated)
		.txswing5             (),                                                         //         (terminated)
		.txswing6             (),                                                         //         (terminated)
		.txswing7             (),                                                         //         (terminated)
		.txmargin4            (),                                                         //         (terminated)
		.txmargin5            (),                                                         //         (terminated)
		.txmargin6            (),                                                         //         (terminated)
		.txmargin7            (),                                                         //         (terminated)
		.txdeemph4            (),                                                         //         (terminated)
		.txdeemph5            (),                                                         //         (terminated)
		.txdeemph6            (),                                                         //         (terminated)
		.txdeemph7            (),                                                         //         (terminated)
		.phystatus4           (1'b0),                                                     //         (terminated)
		.phystatus5           (1'b0),                                                     //         (terminated)
		.phystatus6           (1'b0),                                                     //         (terminated)
		.phystatus7           (1'b0),                                                     //         (terminated)
		.rxdata4              (8'b00000000),                                              //         (terminated)
		.rxdata5              (8'b00000000),                                              //         (terminated)
		.rxdata6              (8'b00000000),                                              //         (terminated)
		.rxdata7              (8'b00000000),                                              //         (terminated)
		.rxdatak4             (1'b0),                                                     //         (terminated)
		.rxdatak5             (1'b0),                                                     //         (terminated)
		.rxdatak6             (1'b0),                                                     //         (terminated)
		.rxdatak7             (1'b0),                                                     //         (terminated)
		.rxelecidle4          (1'b0),                                                     //         (terminated)
		.rxelecidle5          (1'b0),                                                     //         (terminated)
		.rxelecidle6          (1'b0),                                                     //         (terminated)
		.rxelecidle7          (1'b0),                                                     //         (terminated)
		.rxstatus4            (3'b000),                                                   //         (terminated)
		.rxstatus5            (3'b000),                                                   //         (terminated)
		.rxstatus6            (3'b000),                                                   //         (terminated)
		.rxstatus7            (3'b000),                                                   //         (terminated)
		.rxvalid4             (1'b0),                                                     //         (terminated)
		.rxvalid5             (1'b0),                                                     //         (terminated)
		.rxvalid6             (1'b0),                                                     //         (terminated)
		.rxvalid7             (1'b0),                                                     //         (terminated)
		.rxdataskip0          (1'b0),                                                     //         (terminated)
		.rxdataskip1          (1'b0),                                                     //         (terminated)
		.rxdataskip2          (1'b0),                                                     //         (terminated)
		.rxdataskip3          (1'b0),                                                     //         (terminated)
		.rxdataskip4          (1'b0),                                                     //         (terminated)
		.rxdataskip5          (1'b0),                                                     //         (terminated)
		.rxdataskip6          (1'b0),                                                     //         (terminated)
		.rxdataskip7          (1'b0),                                                     //         (terminated)
		.rxblkst0             (1'b0),                                                     //         (terminated)
		.rxblkst1             (1'b0),                                                     //         (terminated)
		.rxblkst2             (1'b0),                                                     //         (terminated)
		.rxblkst3             (1'b0),                                                     //         (terminated)
		.rxblkst4             (1'b0),                                                     //         (terminated)
		.rxblkst5             (1'b0),                                                     //         (terminated)
		.rxblkst6             (1'b0),                                                     //         (terminated)
		.rxblkst7             (1'b0),                                                     //         (terminated)
		.rxsynchd0            (2'b00),                                                    //         (terminated)
		.rxsynchd1            (2'b00),                                                    //         (terminated)
		.rxsynchd2            (2'b00),                                                    //         (terminated)
		.rxsynchd3            (2'b00),                                                    //         (terminated)
		.rxsynchd4            (2'b00),                                                    //         (terminated)
		.rxsynchd5            (2'b00),                                                    //         (terminated)
		.rxsynchd6            (2'b00),                                                    //         (terminated)
		.rxsynchd7            (2'b00),                                                    //         (terminated)
		.rxfreqlocked0        (1'b0),                                                     //         (terminated)
		.rxfreqlocked1        (1'b0),                                                     //         (terminated)
		.rxfreqlocked2        (1'b0),                                                     //         (terminated)
		.rxfreqlocked3        (1'b0),                                                     //         (terminated)
		.rxfreqlocked4        (1'b0),                                                     //         (terminated)
		.rxfreqlocked5        (1'b0),                                                     //         (terminated)
		.rxfreqlocked6        (1'b0),                                                     //         (terminated)
		.rxfreqlocked7        (1'b0),                                                     //         (terminated)
		.currentcoeff0        (),                                                         //         (terminated)
		.currentcoeff1        (),                                                         //         (terminated)
		.currentcoeff2        (),                                                         //         (terminated)
		.currentcoeff3        (),                                                         //         (terminated)
		.currentcoeff4        (),                                                         //         (terminated)
		.currentcoeff5        (),                                                         //         (terminated)
		.currentcoeff6        (),                                                         //         (terminated)
		.currentcoeff7        (),                                                         //         (terminated)
		.currentrxpreset0     (),                                                         //         (terminated)
		.currentrxpreset1     (),                                                         //         (terminated)
		.currentrxpreset2     (),                                                         //         (terminated)
		.currentrxpreset3     (),                                                         //         (terminated)
		.currentrxpreset4     (),                                                         //         (terminated)
		.currentrxpreset5     (),                                                         //         (terminated)
		.currentrxpreset6     (),                                                         //         (terminated)
		.currentrxpreset7     (),                                                         //         (terminated)
		.txsynchd0            (),                                                         //         (terminated)
		.txsynchd1            (),                                                         //         (terminated)
		.txsynchd2            (),                                                         //         (terminated)
		.txsynchd3            (),                                                         //         (terminated)
		.txsynchd4            (),                                                         //         (terminated)
		.txsynchd5            (),                                                         //         (terminated)
		.txsynchd6            (),                                                         //         (terminated)
		.txsynchd7            (),                                                         //         (terminated)
		.txblkst0             (),                                                         //         (terminated)
		.txblkst1             (),                                                         //         (terminated)
		.txblkst2             (),                                                         //         (terminated)
		.txblkst3             (),                                                         //         (terminated)
		.txblkst4             (),                                                         //         (terminated)
		.txblkst5             (),                                                         //         (terminated)
		.txblkst6             (),                                                         //         (terminated)
		.txblkst7             ()                                                          //         (terminated)
	);

	pcie_cv_qsys_mm_interconnect_0 mm_interconnect_0 (
		.pcie_cv_hip_avmm_0_coreclkout_clk                                        (pcie_cv_hip_avmm_0_coreclkout_clk),                //                                      pcie_cv_hip_avmm_0_coreclkout.clk
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),               //                      onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.pcie_cv_hip_avmm_0_Rxm_BAR0_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),               // pcie_cv_hip_avmm_0_Rxm_BAR0_translator_reset_reset_bridge_in_reset.reset
		.pcie_cv_hip_avmm_0_Rxm_BAR0_address                                      (pcie_cv_hip_avmm_0_rxm_bar0_address),              //                                        pcie_cv_hip_avmm_0_Rxm_BAR0.address
		.pcie_cv_hip_avmm_0_Rxm_BAR0_waitrequest                                  (pcie_cv_hip_avmm_0_rxm_bar0_waitrequest),          //                                                                   .waitrequest
		.pcie_cv_hip_avmm_0_Rxm_BAR0_burstcount                                   (pcie_cv_hip_avmm_0_rxm_bar0_burstcount),           //                                                                   .burstcount
		.pcie_cv_hip_avmm_0_Rxm_BAR0_byteenable                                   (pcie_cv_hip_avmm_0_rxm_bar0_byteenable),           //                                                                   .byteenable
		.pcie_cv_hip_avmm_0_Rxm_BAR0_read                                         (pcie_cv_hip_avmm_0_rxm_bar0_read),                 //                                                                   .read
		.pcie_cv_hip_avmm_0_Rxm_BAR0_readdata                                     (pcie_cv_hip_avmm_0_rxm_bar0_readdata),             //                                                                   .readdata
		.pcie_cv_hip_avmm_0_Rxm_BAR0_readdatavalid                                (pcie_cv_hip_avmm_0_rxm_bar0_readdatavalid),        //                                                                   .readdatavalid
		.pcie_cv_hip_avmm_0_Rxm_BAR0_write                                        (pcie_cv_hip_avmm_0_rxm_bar0_write),                //                                                                   .write
		.pcie_cv_hip_avmm_0_Rxm_BAR0_writedata                                    (pcie_cv_hip_avmm_0_rxm_bar0_writedata),            //                                                                   .writedata
		.onchip_memory2_0_s1_address                                              (mm_interconnect_0_onchip_memory2_0_s1_address),    //                                                onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                                (mm_interconnect_0_onchip_memory2_0_s1_write),      //                                                                   .write
		.onchip_memory2_0_s1_readdata                                             (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //                                                                   .readdata
		.onchip_memory2_0_s1_writedata                                            (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //                                                                   .writedata
		.onchip_memory2_0_s1_byteenable                                           (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //                                                                   .byteenable
		.onchip_memory2_0_s1_chipselect                                           (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //                                                                   .chipselect
		.onchip_memory2_0_s1_clken                                                (mm_interconnect_0_onchip_memory2_0_s1_clken)       //                                                                   .clken
	);

	pcie_cv_qsys_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                                            (clk_clk),                                                         //                                                          clk_0_clk.clk
		.pcie_cv_hip_avmm_0_coreclkout_clk                                        (pcie_cv_hip_avmm_0_coreclkout_clk),                               //                                      pcie_cv_hip_avmm_0_coreclkout.clk
		.alt_xcvr_reconfig_0_mgmt_rst_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                  //           alt_xcvr_reconfig_0_mgmt_rst_reset_reset_bridge_in_reset.reset
		.pcie_cv_hip_avmm_0_Rxm_BAR2_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                              // pcie_cv_hip_avmm_0_Rxm_BAR2_translator_reset_reset_bridge_in_reset.reset
		.pcie_cv_hip_avmm_0_Rxm_BAR2_address                                      (pcie_cv_hip_avmm_0_rxm_bar2_address),                             //                                        pcie_cv_hip_avmm_0_Rxm_BAR2.address
		.pcie_cv_hip_avmm_0_Rxm_BAR2_waitrequest                                  (pcie_cv_hip_avmm_0_rxm_bar2_waitrequest),                         //                                                                   .waitrequest
		.pcie_cv_hip_avmm_0_Rxm_BAR2_burstcount                                   (pcie_cv_hip_avmm_0_rxm_bar2_burstcount),                          //                                                                   .burstcount
		.pcie_cv_hip_avmm_0_Rxm_BAR2_byteenable                                   (pcie_cv_hip_avmm_0_rxm_bar2_byteenable),                          //                                                                   .byteenable
		.pcie_cv_hip_avmm_0_Rxm_BAR2_read                                         (pcie_cv_hip_avmm_0_rxm_bar2_read),                                //                                                                   .read
		.pcie_cv_hip_avmm_0_Rxm_BAR2_readdata                                     (pcie_cv_hip_avmm_0_rxm_bar2_readdata),                            //                                                                   .readdata
		.pcie_cv_hip_avmm_0_Rxm_BAR2_readdatavalid                                (pcie_cv_hip_avmm_0_rxm_bar2_readdatavalid),                       //                                                                   .readdatavalid
		.pcie_cv_hip_avmm_0_Rxm_BAR2_write                                        (pcie_cv_hip_avmm_0_rxm_bar2_write),                               //                                                                   .write
		.pcie_cv_hip_avmm_0_Rxm_BAR2_writedata                                    (pcie_cv_hip_avmm_0_rxm_bar2_writedata),                           //                                                                   .writedata
		.alt_xcvr_reconfig_0_reconfig_mgmt_address                                (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_address),     //                                  alt_xcvr_reconfig_0_reconfig_mgmt.address
		.alt_xcvr_reconfig_0_reconfig_mgmt_write                                  (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_write),       //                                                                   .write
		.alt_xcvr_reconfig_0_reconfig_mgmt_read                                   (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_read),        //                                                                   .read
		.alt_xcvr_reconfig_0_reconfig_mgmt_readdata                               (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_readdata),    //                                                                   .readdata
		.alt_xcvr_reconfig_0_reconfig_mgmt_writedata                              (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_writedata),   //                                                                   .writedata
		.alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest                            (mm_interconnect_1_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest)  //                                                                   .waitrequest
	);

	pcie_cv_qsys_mm_interconnect_2 mm_interconnect_2 (
		.pcie_cv_hip_avmm_0_coreclkout_clk                                        (pcie_cv_hip_avmm_0_coreclkout_clk),                    //                                      pcie_cv_hip_avmm_0_coreclkout.clk
		.pcie_cv_hip_avmm_0_Rxm_BAR4_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                   // pcie_cv_hip_avmm_0_Rxm_BAR4_translator_reset_reset_bridge_in_reset.reset
		.pcie_cv_hip_avmm_0_Rxm_BAR4_address                                      (pcie_cv_hip_avmm_0_rxm_bar4_address),                  //                                        pcie_cv_hip_avmm_0_Rxm_BAR4.address
		.pcie_cv_hip_avmm_0_Rxm_BAR4_waitrequest                                  (pcie_cv_hip_avmm_0_rxm_bar4_waitrequest),              //                                                                   .waitrequest
		.pcie_cv_hip_avmm_0_Rxm_BAR4_burstcount                                   (pcie_cv_hip_avmm_0_rxm_bar4_burstcount),               //                                                                   .burstcount
		.pcie_cv_hip_avmm_0_Rxm_BAR4_byteenable                                   (pcie_cv_hip_avmm_0_rxm_bar4_byteenable),               //                                                                   .byteenable
		.pcie_cv_hip_avmm_0_Rxm_BAR4_read                                         (pcie_cv_hip_avmm_0_rxm_bar4_read),                     //                                                                   .read
		.pcie_cv_hip_avmm_0_Rxm_BAR4_readdata                                     (pcie_cv_hip_avmm_0_rxm_bar4_readdata),                 //                                                                   .readdata
		.pcie_cv_hip_avmm_0_Rxm_BAR4_readdatavalid                                (pcie_cv_hip_avmm_0_rxm_bar4_readdatavalid),            //                                                                   .readdatavalid
		.pcie_cv_hip_avmm_0_Rxm_BAR4_write                                        (pcie_cv_hip_avmm_0_rxm_bar4_write),                    //                                                                   .write
		.pcie_cv_hip_avmm_0_Rxm_BAR4_writedata                                    (pcie_cv_hip_avmm_0_rxm_bar4_writedata),                //                                                                   .writedata
		.pcie_cv_hip_avmm_0_Cra_address                                           (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_address),     //                                             pcie_cv_hip_avmm_0_Cra.address
		.pcie_cv_hip_avmm_0_Cra_write                                             (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_write),       //                                                                   .write
		.pcie_cv_hip_avmm_0_Cra_read                                              (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_read),        //                                                                   .read
		.pcie_cv_hip_avmm_0_Cra_readdata                                          (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_readdata),    //                                                                   .readdata
		.pcie_cv_hip_avmm_0_Cra_writedata                                         (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_writedata),   //                                                                   .writedata
		.pcie_cv_hip_avmm_0_Cra_byteenable                                        (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_byteenable),  //                                                                   .byteenable
		.pcie_cv_hip_avmm_0_Cra_waitrequest                                       (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_waitrequest), //                                                                   .waitrequest
		.pcie_cv_hip_avmm_0_Cra_chipselect                                        (mm_interconnect_2_pcie_cv_hip_avmm_0_cra_chipselect)   //                                                                   .chipselect
	);

	pcie_cv_qsys_irq_mapper irq_mapper (
		.clk           (pcie_cv_hip_avmm_0_coreclkout_clk),  //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (pcie_cv_hip_avmm_0_rxmirq_irq)       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pcie_cv_hip_avmm_0_coreclkout_clk),      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~pcie_cv_hip_avmm_0_nreset_status_reset_n), // reset_in0.reset
		.clk            (pcie_cv_hip_avmm_0_coreclkout_clk),         //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),        // reset_out.reset
		.reset_req      (),                                          // (terminated)
		.reset_req_in0  (1'b0),                                      // (terminated)
		.reset_in1      (1'b0),                                      // (terminated)
		.reset_req_in1  (1'b0),                                      // (terminated)
		.reset_in2      (1'b0),                                      // (terminated)
		.reset_req_in2  (1'b0),                                      // (terminated)
		.reset_in3      (1'b0),                                      // (terminated)
		.reset_req_in3  (1'b0),                                      // (terminated)
		.reset_in4      (1'b0),                                      // (terminated)
		.reset_req_in4  (1'b0),                                      // (terminated)
		.reset_in5      (1'b0),                                      // (terminated)
		.reset_req_in5  (1'b0),                                      // (terminated)
		.reset_in6      (1'b0),                                      // (terminated)
		.reset_req_in6  (1'b0),                                      // (terminated)
		.reset_in7      (1'b0),                                      // (terminated)
		.reset_req_in7  (1'b0),                                      // (terminated)
		.reset_in8      (1'b0),                                      // (terminated)
		.reset_req_in8  (1'b0),                                      // (terminated)
		.reset_in9      (1'b0),                                      // (terminated)
		.reset_req_in9  (1'b0),                                      // (terminated)
		.reset_in10     (1'b0),                                      // (terminated)
		.reset_req_in10 (1'b0),                                      // (terminated)
		.reset_in11     (1'b0),                                      // (terminated)
		.reset_req_in11 (1'b0),                                      // (terminated)
		.reset_in12     (1'b0),                                      // (terminated)
		.reset_req_in12 (1'b0),                                      // (terminated)
		.reset_in13     (1'b0),                                      // (terminated)
		.reset_req_in13 (1'b0),                                      // (terminated)
		.reset_in14     (1'b0),                                      // (terminated)
		.reset_req_in14 (1'b0),                                      // (terminated)
		.reset_in15     (1'b0),                                      // (terminated)
		.reset_req_in15 (1'b0)                                       // (terminated)
	);

endmodule
