// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:05 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TyTSKKfvj8zkI9TVgYSNdHgI675nlmgKTRlb6WJNaH7379MGkK8FFBo7dS5eNjMF
XK0ZflmAPgr+zhGjAeJjdWk4Uk0V0Ur+mvWxiB+eTNB6fvoywzrJqszKeZ2y/TEN
1WYtZUe/CuStOhkxyOe3ctzogTvKtSwogpTO3OGceSM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8256)
BiINaewamgZRhRGJXR7gQD6Hxqv2tVAaQ/GMVYRxGniq8G6WJXtB0EK5KV5qqcR1
b4JjQhB7ROem8LyxGM9iMe46OZdSnAnoQu7bhsM58xmqlgV2UjBJecBAyUWtQWDa
ho3kcx7acdjLGrPR/An6jRSNIfeEhU8a1tP7xHKaKbB6QMLW9kmkc1aPcdRo/P5n
23o5U1Se/IgdxcTwBdX4QfHw/+qaq9xBmfVywUGeaiqIm4kYCb5VKe0iXsU2KE8C
XAFCLDQ6kfIXR+H4hK3oGo5s9EF8ZwwgSQRm7d22czaTGOsXdY4HrTjzrb2C3pCg
SQ77ZgbYaf1Wevt//eIuFo1I4S+66Bc8lSwlYfhIPA8zZXzVb2kbDhdIVbFl9HVa
9EGrfP8RLlVw7vp9tMJmvZ/8dHvz34iRCK4yvX1HC/4eJpKKjtqVjB9SuWp2FBQf
IpJiV4T1S9Tjdg2V9089VQaiikZCgDfKLwQ+poOI9ZtnCN0PN0TuJKraAHAdASzY
vRGNU54KHX+PBVf7c0UHoEm/ouNAUfYIm7F4a6NqeVWsEp4VBLIE+lTV9KcW9+pn
5sBDyyhCi8LvmdH3zNt9UBFELVeWxuymUvmgZrZclx2N4CnxDEKrlYvLoe23mfSV
gCBMD6EBcPD+rcfGMyHAp00eUTpFdouLOenKoNT1dBMq9sbqlqLlfstWxBtoTGzV
bykepNlBlHIRCgnxkP/cD/ExqBP0uFzRTdqiIevsZU/d/FlIJGJvw4ZkqvKeMFc+
lKdbP9qU8aWVr90376dT4JH32GI3D/QgJ+iHphffBz4VjvQCb5tuVR0arhiTOBTq
jJNEyDOVfgVhqOSAjXtam1vBNBly1ZGEpZ9rhEv4LLKg/nXo8nxS9n6YnRJBDp3k
dJ99MKlT3v69T3zrAzK5F1aZ6z1Fff40Ik7nHdpBPcYO4v6DE18Fw46gB0GRffwf
SicaTDfNawqcr7+xBudhbx5fuzYzZ8VhqjFhw1/j80L20jouzIfTPF3mWdW0ZSu0
VjyN90Z/VuPoSnzwqhf5r8Z2pTuaKA/Rk8x+sK/n9nuvHA9X8c6DyWTnQcrexUeo
Y3a3ysqqg0+SrIMqi/g7wxORrF44DGqaMJoIPDLu2TolAJZ1AlBufFDlh8Jd3Obz
YkUQuQIB9Jo1lph3aXWnOB74nNFETP4QuCGYFdyAzgDXDdeqZ/ACK78esrg5bwGH
6hzwADG2ZGWiA0omIFB1FUPHI66WSBd5bI9K5oHtNsRa3nBuyFzAhWJv/+ICWxWh
83yS1GNH0bBsIaP61oYoX7x4/eN9TjgzsCnWXi7B27TH+TZdazrO9PDaCm6dm9Jz
fLVE7mRd/WFLgL/CalrhyNTWaEhpPs5nOT6xvvIyzQQLaVw/TdtdFbA8wuYcPCoh
0b602njbJk48PXOMY+Ip7FJRWa/wquczWaRQqDvPe/iCfgxJVIJkOpREJLpt2P4z
dBWy89GQOEe9GtuUSgp4H/E5F3Fj09/usxXvVkSrXfy4nKZdHvbyTQr8PXOuACph
dtJao4edV6+R8ReKNYRwqQxT7EBYRxaCLuJ1/Qjp3jxQ3/WntOks8i0aAIAHZb5c
ib6SqOq+nIALsfy7oaOkk1nI31LPawdNld/5fKrIVi5ztsop+Z6mQp05CuZXMF2i
IkKolUctKtoqL3DNKYxsZR6sZDf0HAfTwdOmVosAfzcYwBG2N3bR7yCmx0xwvEob
aycUIcyQ2SUHPLLgC9BeC+689p/4cil5PAvVY4vCm+OkRc7I4YscYeY2Xhsy5W+X
BDoOSn9SpmYBf6XbzzUEpY25vygH+71IGXZzjQk7pluRwMRS9n7HrFceUpRJrvwz
NxERxPUOAdUJVmDOva/uLwjRxlkmPWMbHLQJN7XT/yX4m8MG22tR9RqPjbdZJyew
souLwOOp/mkkh/p16gJtmP9b6DLUzOOc+szyf2U1cL0KmhYX91hHuNPKYlRYqyaG
GAzB2vaiBtM+9IytLYTVpPk7JjruMGXi+mo607zVoTSOpDgVTlO0oLz8Xmq53smo
oGRqu1S6xrITWg8H0hc0SWQY3O6i9TBVRjJ/rsU29tI0zJ7frD8cuo62MsSDQAxV
S8sWwiDITUnnyYYF4wza2NherWV3ThIN6Bda4xRztGHQNEV90swsZRB5MBRoQvwf
QTItKbIpRctSqy7SqbMPCOqBRhZ0/tm5Mlw9KbGFe000IoIcaxR/OLucB6Mq+Zvv
jbNdEWY89UfZmAIE/TG7NgROpb/i/dLDGF8OYehOOyWpoK6L+zXMGwoGgVdtQUQh
Fu8G7NT417v1VOV8wXUw2EIhrtAiXRMmSQKn0r2dcrGZOgHzREYcilkhDOWlQ5he
m5WwOascw6l4yb85Gye/olkfUEs6twlrvfUff3Pv4mP+RgaYrjfA4btTg2pFjbIT
PWouIpZnKv9fed1qDPG19qimZ3tP4Qehle5s0CukrPl0SC7c0fTGspchqD26INry
IWKjAg97dMwkFfFSJCJPm6iCqvd6p3sDkugRtF4VOQq1wApnb+Gn+Ymk1LYJrpP4
4m5CS7yc4gZFNcauGsFF3Kj0K8mWWF7x6tFYPa0qz+5H3/7CEipMRVw5wK+X7I/3
TC7PAg6TfS8gOOJoa8b4sNNAuLgS0wx41bowh68zPLAwWyGb5q3aR1wJ0xpaqMtR
yBfXHEtj3ofjWq8H6r/wFp2OhQWqRdtwh1LcMJ3qLcBT7Bmc2cZjTyyi83lEcV3A
dvI8PfLpWquDYBNKZy8DUc/7r33xb1pHxKrIPEH0sAyM/7OWa0JqJp/gxO7EiYfV
nI2RLWmezHa5piwYH8SB1jgqMEGpqRkejFUw8xWzjpJ2VJjmvgqJ2fdsaFLaR/HG
+Y6Ey8aVXyn6Udxnbzg+PLN7s44Mv182JQyCZh8mh4s/my96AXnvCtKXiYosh8ki
XITPRfrb0p3Ua14qAvjaj3X7wyBj0U9q2TX5HdIwqrw4PZ64qAsdIA0uu+GuWH7m
zej/EbewUAGXrrfxBrtzGKZ/mtm3HleoFatcajd3qFtQd6+fyosJfmdhDAgGd0Qr
rJTmSexwd3LkQfcLuNlk4gUlMlx0L0W6ABQg/xc20DkwwOQ1s8cNquAdH9qVznhn
/NY9piPZOJHWkKjKPL/o7N65n+aBpUfkwVy3YYre4KgIkZCZQzVwNutAV16nMPU8
3Rb3+Sf+Ym3WLxMGiXYZmI2s2hqi9ddv7/qauReb7BqAPTDAC8kAtbucnm8QFoKj
bXeb4hTHaXU36l7E2lShnsb+quKe9rtDI5dkvxiiIW28pgjC+P4dtUHD/cd0idV8
QtH8yJFT4udR7TiBzGGRLkqdTGer8xeDOGKM73Orh/ES5jKz48udH4AsnaZ7e/4V
l7I/AGXNoP93lajKdaq4fwCkj/NK6EbIitdO+KV38Ci0bhRu6bKxxt4b5fSQcDS4
YPupP20lRBUsQ357qA/yafPfKzWZDPL33FP/vdrx88luOmEzmm638oNQoXPbfNyL
yz6jJmne46ZKgF/J0dTstvFF6P9JKJHZwkEBfd7RZ5VXIN6fcslixkJbpsZsq680
nIm+TyeN/vGQVvb15cKcVjogNJRa95kKcbs0CK8Oafz8//EnjmCkyNYAVIf8U0qp
oaw7rut47Xv/yaxKIvTZhW39ouzcv5JJjS/4sOKxasgGn/gGaO6GpOAoAj9EDuwD
TU7mJawd27GFYkIeMxOP633ZOwzj2zlRlw0YJKgSUdLJ7+FU2tXQ7t1A/R3BqJ+Q
a/TiluU6vq2WGSQ4P2zlon0wrBhK5j8q/9NRGtw88MqDW8/B02RprkQAIy95kqdS
4eWMhF63INvu+Ts7X4QKgskWCc9GMZ+cVkBNqiXKt+ynomHdCV3X86LLPqW0geKc
I2fyPcd/+ouacypwNwrkyvgkEnJxvVamJc710qVqlIRIbFd0J4DIWdVC0AqBNbRa
QuDR6Aa68NVELerHYIbDHSxzZ3Bh2iSS5XXgmDLJs14Ef2n6scOVeb+oqtp+PW/k
nCOxEXNcf9crHLLdqlSPjLKCzpsFrr5Nd4PRAv/eSPO9Io/y0/XqnNY8HXAcztoj
Ef18MAhEqBWqak0WHBemUcUjPmIkNrE7GXwbPjScraoacPWYP1gfIq1UO02a18c6
RRepQLbqZOmnjrWg6Lz6M8XYLPIneHnOVigfTJjAvZUiX2vC64NWwQSvSCZgVDDI
wFe6cEpZVanKTEn7H1Cd8/PqqpgW+/9Q+fgzJQ08ItaKw2NmNCvMRA9/OUyCGk2x
CdMbhwmJCLOc4dhLG4TThopMj1XPXmAkgF8dxNeBcoPY6WZ/zGdc/mTF1wHEaf7F
/yCM9jcWq3VbRJe3GXSZsBsML9vCOU8RqJOXrOnNnWhqK6xHEq+2dEJ0dmilQMcT
y3gSl7DmcmJVDfrugkO4K7cvOLEPcayBFFPmWfKL+qIGSRFbfRLgbzDaSMK89jGo
71Q81bj9+ylvDJuEmmuI9roJ2xKnDpYOYgmlymcmIp/5IfF4TlyB9zD+IptNoNpl
aTtHqlmWEpRtdY++BgvF3VpOCFN2+cYHqC3cPVlep1IwKJUdpQOz+4I5miYVztCJ
E4oOSRZNtYQxD3sYLT6M8SnKlTIcV/oapDiB9bz4XHIOJsZfGiaHiwMpjAr4jwuY
XaGwRsSSeEuNjWo7jH2hjJX56aBxkNpbU6sN1YbvmDWBCjlL435QQsptMeyrNQW/
oXHw15AzroIzqe92zWvuM1wKRZLYEHUuVo9VyonmoCwibla5FO7Tuy/lvVpT9in6
OmgiMdvz3cICOMxcWrpksK3afSlmuS5Z6uF+KdMrclgCnLYBuaGXJnhdSkyndsO7
lutirwJZJS3N+Ywxtw8WkQS4u3nrKYzS3e/zpuCWruSXK2+63uS+4pOgObPD3ZxB
k2QhzpO24Qfi8QEr7f4cKk3TsmKhGXsOe8Cii0PdLXixHMF7/xg9+ehqnNz9VaI1
jo2Ui1XzC3kAjHN8dhTxuLtcpHwvTjjeD51N6xbMkGMvM4Hm2cl3ESoWEYZvgOWm
MF/sJjmVyNWFDqXmq7A5ciqZCkwwxDHTr4PPu2br19ZlTycRNJZhqap6KrF1lhxR
Nt9dqKjDISi5vx3CLcXOdCMxDzoOUqh5v9bQn4kkhEth9fFSo1tB9bn/KrprS8Xx
KpZE8cwDVs+id8/T/pGQ6owvpjEq+yj6UUANQK/Bhb3kBgsTVks3vaR3FLC/bfl3
BpGLGIiJe+tjhxVT/6sBVsll/WLIJinnELSTpM0/lDdaGSRlE0FWqV+ZrUWAMvUG
6pZGw4UVSco9QyrRbVjZiRJBIal35AhXjEU9nX1EGRqPSLuyBR9gotyqal6j4YsJ
lK1BOrZ/D0bmLyIiHtQaebQphxQJuxJQe4JAoxEI8guQUSHX6gBuBaLtJ6taNj7P
4exYvLDeGez6uTlmXdXHK+59VpbQ6pt7LEMy+SR+LexTHsMWHiqk+QvYFnJuty4D
E7xcDDJe+eD4Epb1wVld6ZamRzjmPFrsZPldWiXykhnaIhDY6z2E/nVMlHW2S+1f
PcPkKN3z+y3Fj212g271bpv4zzVXU9skPiOQNmHaNJYa8aVRXVvUnqzN8LLZvb+c
VqZ48afSrByDfmMNsz3710W/ixe8x80mfmVkSjDMkbUqQ1uQoHV9DQge5Yi9QVmP
7UfUzNgc4oR6E4bHpfIUo+pn8oa6+d0b6MdnfOmCHzCwUVH9M2KDofGLmtasSCMQ
8hZi+ZcqdrnYavLN42ccIfIF2j2S3GI4w0uW5LjAc0vWWoDzcNfzMVktq0FQ7pLN
EKe0VqRZuEgclcmDB6jitpvvqbw4J9XaADYHsa6PAc6CM1y1XGvNSkl13i8hrNRf
z6NinXy7SbJgZI21gEqYcmRHSFYgzhAA1AdZiqCBLZb73jD4a43ZtnbBWgsPc/Fo
XjFc4t+gw6r60+oKxquCsO1Cd7rOiuvLqY19nLPROnYFXHUb675k05p5r/ux7Qql
blO3Y3NRH7rAhI4lVFjXGQBD6+rb/rDdKzUTNoMu8viHiVR+ZdrhNu171tNkJ1h0
MYCACBRFCb953hfQQhm1BOFSprO2RjXKOrvRTkbQvL/BaL4IPV0f1ZHu7yDMJh5n
+6T76UunLR+k7VuPbXOuCxLcO4PkjWq+Mh1n3pdBqfkPx3365+AVsSnQPNPKnWGt
Hvw3cKKoR/nNYV1A8j6TqEW9Etdla8rPl6BMOwgqiIym3q67+lrZmjFU+Yv5eBdu
T6nASuO6GB4sQSz1OOzIbug5zVCEc4Thp6U1ciYdNMxHDji5Sb/ALRXACZ3jZjEw
n0exioYARTNGVDQxt5s9QmUuBTL7XAX13B8G9cV8SBHlbklty9KlEjj+tpww+cHE
ftbrKBQR36Dql/ndqtkade8jaFoV7ejAgo+DNmnRU+J6H2g6FWSIjPXuLNJv0h8o
v9hKmKN+wP157qYw2DG4hgzMr77WRqP+i5+J0joREg3D6m7tBw/x0fku+MdMrzvt
2hXuu7kElkTQ5Gsqr1xmaW9b/mEikiwA7dW3/y9rOCsGx1k2V8PhFuxYrHlGtyxW
LaklCEJvvPrK9qStjjaag0vRA+6WADRZlG3uPfjNMmwhGXz6EVO7xY3GRV6E1cXO
wWNdxJvBKtocm/4YYCZV633z97b+4IKi0+1R3bKYL3F2qdDTHImkxWe0kRIvvznQ
CbdfP5kOXYFhf6ttkzJdv/q13juKo63ZoZzTyXcaRK9akCrG+I9PnjfuNDsF04w3
RJGGkPDP8HDhmFXRdlkOlDjdBfWgaAahxW39gZFppf+Sur5omCeAUNxfdgyCSZOM
p1ThGgHssDgDupf9rBRoDQNVkQtgwOfwJeecl61rv30IkhwsUKnYEvr9SAAF5bSN
NBpMDd/pl6VDDbhKNHMITKb+JQXgtOBFYsXnMX8dRG4LXY0yrd/n7vnmxzOyc+Uh
BIyJW9TF0atheVk8pyDJawftSmfBzI6dQryCfnaUb6xAdzI1tqnfKKn4huTWy4hq
Vx6GyQChdawk/8ArjVl2mlu0mvSl/c6UQ44hay1D+Pelpa5CBSh/V1CirWAAbpvT
RcKtaNqtBQvaJcAhqFEjLc2zLN666TUV9PQ+5fUKixRErUXvFgScwcrJAKNl8Z1N
viNi/IeJKzPS6lqyaDYQ6ODwP0XmwrujOXxL2uTmN6Tuy9xKFQYd/FjEmYeOzPYQ
HnJge01z+ceuxrx9efLKshvz9qePrY4tRaLZBo0Ytgpa1+3KvC6dYscFoC061r/s
/nphuHUfMp3KgUmOAWNESnGTXZL6tzMeJvR2PlfmszIJ9qbgJ1Ha+8d9SkCHjXzJ
tbIhucYpP55PzDTPesW2bSW+PnuoI8ZahxmDi9QAfgWpMMXy6ljXUQyDZr0zOM+K
/Ubf7nmA0oDdp45+/XbWYQZzGPZQvmp0IpnhGBhzXzqzlx1NKblXMB2aEhlN3WxU
ljTxxOG6Wj7cv0PTXVCOeKt6lcMP+ofkshGaObuXPMMkGODYmy+y12Y3f5uXf/LX
5BhLAAujVFxtdpuWzLgZFg90iJi22npxLSq1mCp9Fc1XBYy5A9QfHXa7SPhtKEEy
Q7/l2KBuexB2VCjCZpmy0FH/tpkxUivk4v/NAbM5zjiDekvZeNz+upN2nuZLuB0a
+LZNKf4cbkvWLMgCRBgW/H/XCTdcH2sCPqHLKgzw6hOFys/xoucczcrW63JZ70iK
vklDTVUNYCxvl/abB5gN6BZfXQVa2UE8FcB2znQZvFR4UoDTiFvh07WXVFVAc8Y1
6tkhA2IxoIYf8jRH4rr9po9zVdOdZgodzSH5Jgl+R9WSyumBN/YPvXBLmyfeThpW
O4dnOJiV5JNqJgcoYSpVdpI9tQCqkMRdLwrXCb57l8ugPl070aFYfiG2jHOihPbS
wZx3Gdx3PHErzc7yAegUkropXNCEXbZH7re9VVmtSE/jPQL6LE6VrMbg/u94oIyk
nmy8BxpKc9WfciWUz/swT0HEzX7aedZO3FHOhmW3JWd9fP5It3OqFIWhPoEoIrOI
WnLbN3T6aekMYTBo015TEEVqViWm4cT/X4qXIbhkYB7nFNulybT5LiflOq57/f+v
DXWHYhj8gr6G4TWtVhBpjM3Hwm8QHlllKcrq9dYJgU3nnfFAh/GYJdvblkuqGj9v
uYw7pdxSwQ6PaYHf1EcY3w+kKvPps2+UO5wFyaO0yTG2mQQhUOxdb6BV98D3bvG1
3bN/8T4gNC6z4jeirMZEl3a8lPfxf89eRlAzwN5+s0Upd+uQUkaee93ljDNd6acd
M3aUP4AiiJx4x/zZUoyJJVyrpNNUNaLqWjAnGsY3hhyz5thh3sRpoFuU1FW1S/0z
9NYs3NSlgV5p2IUGdLGpxJJdgONweI8E/9M6WWjlnS700/rTVc+liUuNkhtLx2sk
gNHgu0jpMY2i8Wwg4O7fqMIJ6XYlyRgMyyDwIvTHGPoHb5HELTEuPucO0FaW9sCY
nRvKARljrYTCys6yvbFRxQjB39dpxxKglub7W5/l4ccFGDWfPjWtdS+mm6xnNpfb
hyVBgIL/OI3R1hYm0Vj89jNAHE6rTsDeOOFNwvr6DrUFZir1UIu69EDTYEI+GLYy
pehMNWAI3kOzMTpjADYW4CSSDkJIF0188RDa2cbVggD2PImNC5Ab6GNAsbxHjC50
wWqyKqLM4rB8X89IEEiuL5gmiyE6UO0DXxwaG4ouE8Pa7BDbV4deoMd1hc5UnEU9
avZTkL5YPv9xadVXcK6ImsY8JDLJHTvfrhAD269oLeUV9Izzcyhb/P+5o3LpThdM
bb1GaMRJaZpTyUyyM1AJPkbffS+EIIw4vs+ORZkbVwbtXmJrxJQ6Q3bS7w9+7Jhg
5Qf19aq5fBfKxCyTapveZK8JqQx08X6Aw0cOyN9dMmVvSG/Imyfki+t7lS4ItDw0
pLyu20GFC7XD4VAQ3dLkMiPwSg0Nw+wjPYBxWyDIDfo0r90xj8Nkh4preqfcNRv6
Lf37a58uBdROg9uhPU5s07KnzkRSZDTXeZNV9hoJNVuTEi+aP4/pdu9JG07v+q51
egm9WoVnT74U4vUNhz0Am5XsGZSnEi+j71vcpJftDXpKSE2CrUJI5nfGUYHvSWNw
SNz/o7u86ML4xoXFtnZK/R5HUPSVlWxjrL8FHoEymEXugGFZwnj9vggpzZj7sGcQ
ofskth2zGQc+IHQXpj3EdUGvGuBXGaF5mBgVa/TxE0uUm4zKGVzRFK8vcKsGZ/98
VKyGILc7+oNOVb4+G8mVB1yyBEkq2LFwbmguV1dEpgWhc1w6qFiaHrFwHNDRx4B/
KskWB3DjOfPt3mWIhsAAuDMI3inWh8buEXt4g+Fp1kJ75V1v1T7/wpeV1LDYACCH
A3hUSU/aFPwBmcwXBGdiiE0hQe+aDi12RRxFy2btavFc4mS80lWoTIslg5RczXAi
1Vs6XdgKvNtKJqa9ipVnkduZoLWaZ7bvgMw2qBRRysP/SnaBOMgQK6PlTvKvsFkZ
dQe9xPczUBW4A87k0lZbleRQzd2J6yWqhrxYroatrJB3MP0zxIjFMUoZ9iOZvbJ3
iR49JWO/2ALJvctvgTir0X/OIzFxceCkFzAFMEgVNLtSRseuvVKEKM5+SfNp3S36
5R3PU0docPBG/n4eJB/UMbGRGdnPEgAGVk10ehgJTKusxkvV0fWsJ0TRRS2m6y29
EAClhhojDSlKG23G9AzLJNmLE9ljcSObDoC24JYBl4YsQgXTJFnKjDQggquA24GV
/gGQbhEGKCXGXAOUsWOjBL9aV75uUJaq2QovppzwOk9iO4EIBnoCc1BN2IfSXnza
m6i38XCXG801guibbRVLL3ApGbsRntUbir0Jf9bMPYsllOCDrvzvvSRkXgiMNQeS
HzrRHyBmUEyCQBWhBidaY/tK6lGqS13EmuhSxkJUrZF0Jr4kzeZcqsm3c0S51CSv
htAuSLg9w/e5Elx7YFhmU8FvMIy+fTtMENiiAHXAC75TmfbdVu08F3Ubdtmn09RX
SAPG8aNXZmKktJUWugygruBjtFe0Hc1aWF+CQxdpgKTXh9gJalaQEGR8zzmYsymJ
gkA9fJhYUVULwaUsUESzPwvB6nBzsZwYKrb109yGo3rClGH+ZeG+d87UoxUJJrnu
1arkFCA5NlNOuilue879wqVatd0GSBY+2nGWgt/DXL6PcHhuFktfDTMc7UTVfMo9
qTX+a8HIVMyvZFhXzQ9YTpQkDtDay0JXpTeUV7g/JVx7V7aNzE80nS5dW8+fqwvs
Zk8pnix4qIZNsF1w8cjTv/lVv5jYNfbvCK+JvYor8lJKoyOOxXMpQSJ5N9Jd6pMe
4jQnBJJAfUmToU3oo2fZroscmyt/iKKZvB2NYfivAE+XmUBG36RhtI2X2nf4JC61
JB86jKf18kT45+NFam6U1/uMNH1vfZ99taQroxpMuwBlhec3BJEl6hzIYbFIEUOc
8ZicqQeCvBtCHkTfBZf3TQ1iWhKa+0Mn2UMmE96Z/vUfwYf5smHoub2yX4ITbSs2
YvK0MLG7RBzG9PVQyhg6GCKUQlu76/QARouyIAax8fi86TrLZnH5EE4NPPZeDJWY
gih95nREkQHmt+0JK04GXOxqt3jl4GfDG93eH+eWpcIGjD827r5ABKRhxWdOKsvt
joyFOS9Iv8Jc3Uu+C2FZkAG3B3t+JNV0MXaBtgTiw1uOGJUYhOiUmXxxjYryhGQg
CaeF/UAi/Kp2ZWZHP3K/jIF/UX6PHDi3I1Coco6cunHySA+uijy0VWrubuO5a3OI
nBG9WYDYYbbiSc7+H8738j9XkvL0YLziDQLoqxv1z049daXKPk0VbNzO2Pd3mNVR
M1whixvVpdwIZcUOUPJDOT1GWvinT7LNSx8sDgAT1mPIyCSh5NxLF3gH6/iDiLv5
FlybIs/2y+yEPcsKrwadZDRbzsiMxOAgSGjkZqXKfEEleo/H9oXAH8EXkEZ6zU8U
`pragma protect end_protected
