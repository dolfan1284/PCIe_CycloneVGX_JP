// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:59 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WbMFr6s5Q13n2WWbER/6XC3qsZsBJT0cfvsQUi0aCBocQxswIhliPebbzufXL+pc
eeqaAWYe97rUJyglnloGJpGORNlrItcGPca0GgaB+5Vn4apJpauygxESZ6bqCepd
GEUdX1v5EnRl1kTz26heSx5C+Sg7Amz96RC4fOJX9lE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
CHiHx6esOAMJP6bQri0gfUbFo09xbB27dk1eQzRHSZYEgFJkfZRBn9Mv1ntaE4yg
pME9eAX2a4aKiaaIXyOmb4y9UBlE2uFoH+2Qg5KAKVQqU5Rnlaaq2VauESEVriCO
dgNKaQczXHPHVZmMpJ6Q69fcRXv//LoNZtzKHF5S4pyZDnOWSRKJtLxYkl9iK4l7
NJMMOMafBsxvG15rqMgL18PI7Myiqq7DVs8G7d7vkNBjJCDUKoWe7WOMFqbbPll8
xjGglMFJsmC7lijIrcM2lou+o+8oML64tcrK4yGTET92ExCebOadkSnmXYUR3QwV
kk4yloae8qSc0goomU0QMZj7MDkCKuXiftAfdbmHjPtO+zg4erXeOjflviBS09tc
Uf87CJ2K1/DTflsbSfuoxzo4/Hb47kzx6CaX1ePZqBTE2tFj6pY7e78Tmkt7nd3+
5RSXJWH60qEymiHhoup8WITwXHM+ABtBEMVR5yuJq3zWhuXuKLv5oPxsmBtaKciI
ocI9kWhGA/WD9k5n6K01Kf6mzL2pbQImqH7Wroa7XgBzVVmiJEhYBqJgtvURJuBw
6bQKCiIiAzPoia5lkor399XzJ7NypGbfNfB3dt9V2qdSq1jqik4CxtEKdtlR7DoX
0U0n1WZp56frxdars6gov7w7Fs0fKGJChgilWKe/3B1YpBH++J/nwrN7ahF0J57d
Rx+TfowfHiHrUy92096CuJkwj3Eh01nOwkMopJbqCk2SrbyrUOOS1+q4qsn3lNTq
6MzVtazvg19JSRY9KfD9PGiwQ6BJBxifzm0p2uz1Lm8c9hsSULt3lJ6zSc0F/jLn
IKmkLRdWTMI9Ydt9XHD/2RGDoJpH52vVFVP8p1MmS0IbKS7CQGdB4Yo5XTFUAMqr
crVkADNCjUXeZqIFVPhnD654EVkxA8ZcVF8wcFLEW0YuerunEXipczzpusDd/lb2
eNUKzSYGcPb6Uxf4AXTqh5AS35lAIgXx+rxkEwUuMLwtKPjDIhuLI7PGU/vp7uW/
JAtnjGjp3R7pzc7TlWHFiV9kdSlruj4nALCGky3b5UHKA+QV1L0ZGMoVQnF3osVU
zWLSfvWmXO2KbI/DpAQtlwbrkwvF2T9NPj53qbkKsyuKJaHNbR+whwiOyY7KlSlL
u0EdoIxRipKcU8l5wdDXul1DPhR/JPGYPKVVclbXhjFXF8k7FFdoe2YCY+hwysMD
fi8N28yO4o7kU0sxcMNl746tdeWddF7zzH8Lp0+ITsw5/vjNMWWky3rtpriE5xOO
MytObaMRzsM+T+YOJ2XcICFIbsGGKlnJKPbdv6pCpHJkoIiyy51DLmMznHzES4+Z
NJZvuarkqDi+JJMsdzLh14eFAllQ1Bj/7Za+5liiA3xoeY54YHLoAg56ElyXK3MY
z+6kqs3ddkrEh0kO5wn0cWBZCSERR5YGdZ5uTFwljcSbAEy/1xk7iCQubq/WEkS0
tKfCRFhi5cKtyDv6nTjZQfq51+u5QLn5E11QdkJZetvnGp0MyLRV4zh452ag8DIR
slSWmFyTVKXCKakKLpNMMP5kUtTZI7PBSE0Bmk8kUZxfWvEChnJT/qGHNnEm+Q2N
rapO+ywF/tjjLpbuUEyyJ51I9tDZoGT2wp9KodmX5Z7vO3i0XddOOTWu1jA6+qMG
gkaaeCL3Z6UNrApIv5UFBy046l6g0ttU7YETVNN7UXLj6wfPmI1b11/xNzXm4ht7
FXPSGOMdCqR1y7xsEATV2PFLoIatZE7N8eN6BI9JdiNQ/uZklCt2BbJCTCxjzeg3
adxNf6NlBI9p4eTHoHwcmoAAa1YyaidyIzB9cdTesxHqvzD+vS0A5OxCEb712aiq
0s0v1hJLn64WAkq1CPfvGZW6pb/DJU19S3HAKlVX94wK+Wj+DsByI7VRYVmx02JL
21vB7se9wBHhGGwjL3x1XMUwsGSFYLMnyaWgP4nHcTGkpUdNcTl9JEjR36h3z7xT
fDtMcyMF53HsmaFVkbl3zSODIoOQVL62wZoChD3dbKNgTfWsDotc+kL4NXI1FEqZ
sMnVYOgooObg5yDWYBtWi2+9GtYRZxJ7DJ9Bq1S3ScP/rERFvjk3mDtJWRLLkBoG
KY0IU1rN7+L4zwR7xpC4dyUajpWH6IRdyBhaaRJwnpvWqCZcDtbFiGae7kFJU8WB
NtJ+fIe9eU0IaMfOQhMXML37R+08jQrvRxWJVBg6v126FpClm5IoKyjGRxqf9Lp1
LFGJNAruBM+niLV8wc5bILVJcKNGkJJcs1haYhAhNTEItGBN6PqCIORwGgnOyKQu
gp81pXIxQ2Ulw8CC6FniXJKvHYmIu+SX0iOKzVJB+5EAVQ58A/3KhHLeYDy9Ryah
7iHJk2gzilR3k6jwSS6xgz4TWkmVJRNsoDIBsHfE/mMfPMzPHUf3yDbOUPWnWJIe
ioJAgfYLEoz1cC4GrHCAV8dlC4U0YHx9Mmz67mvCTQa1HhGYTHFABFCc929wSfPm
mYNXczAhBoKQRoWosAH1kZyPgfGxEG59RQwGuv7eH7gZIw/qQKftIiDe/y7XQyuH
SU9Y4x6v6j3iE8jTSvj9F2wZDlaqxWKkbVqUecHySqzps7Ep24PP10nJ4jiLVc5X
Bs5VvBiJ42pCWRrxugT2DSClLFlUOwDPlg6pAiNNfBeiRu7CnEKoHLg/Xr4AdcT4
P/kmep6w2QAcWG9fV3h/KrzUOsStfSMRSikpctYeSJizZ7McoetiWuYpTZQq0w2n
eOya0KDqUDx+seEIydpzo2c7ZJjMYl1PrnoSOWI3ZLy8SqQKlXNRbR0InIyWCmJN
f1fXn9ZFKVf45MvSVBH64s0M1+RAVvRvczQYPd4oIfdev42SbG5PCPan+TnoPJnl
ZHch180waBjs3Dd8jxD4SMOpO3euc+ZwRyrYlNWdUJGvyWA8SxfATc7A5XMYY1xZ
1fqUqEXecCYi0ihYbHDRnrO5nRLvrNCdGg5cVHm7WrJNs4s9+myLrunJrfhcyBG0
VwKRNmCuwMo0zQr18qLkiCWYo1Fk2KZlYMYq4vrCVtIsjpq3IkhldCKg/4xOPUiZ
mbTwsa2w3Za0tbcm8LurSoPfygONASTPFLm/a2HgBgGY5Ahoojbyf+VvpHOtCvi6
64j2b2kleXhPxVH1LXvtudhckM2VTJD74NibwHwRmIZrGhU6ZHR6U+tzHtSHVX7K
RP+I7r/elPAG1aCVMtdLuA7aRB0CNLdFEHWLISy2nFdTyZVKEBHVw1XHu0Y2bVYv
qMPth32r32P0krrJPJWLmQRAHdntSKSAKcCP2/lrHGiBG4yv2pTQypNUc+hyUxQL
KYeYscyw80swrS4QY7gV9d3rRA/JCETBTFD5zSwNXpXLcYMiJNk6mnX59VoUKio0
4bgHksIeYu4tWXzCPcQH38I+HW/VPjoY35POPwLAA6Y0LuZ56U10PL/1wa0kSFZG
KSEQ0yS1HNyC384Q8wPQiQuTXkUNbSkv6yFBVZ1ckcmX83omQ6HyRDPn6CvIwX6g
KEOLPIvbQN9KxaedajkDJmQRaDJtk929uGRqMDsJPrH0hC29fLaDytkDb1MaTXTp
431H8HLIf9JsRRkOjAkXGpyj+zT7wUDdh57mnEjQyWnsA8TPn0XP76EiRCKQ2YAx
trTFLz9Dba3niRuzEoLHIpIANadwTYvuX8RmEMM30Ucn62FJv+6JBISatsvPnf3F
0qOUgNKIXY9vOMox/PNEQY+kjHPYpINwfwGwYOTSryc3q2R1G3r9uECN9SOhiVOb
GzSK9NiOFk/BcaPvTATl1r015dbkUOekQ+c9vfbYhwFz5SKjTOHUiaw6127C06aE
P1VHW9NnDnRAs67dQlgzZsjv+DKLHVjd4RuHoFpMlrE2KsVQlONZBGuKKpCgVySo
u3T/wlabX5ww/IO/zFBmc0PARuX8B+c/P7DaWJ+VL2+M0hI3UUa/a+81gC77JeWg
WP3p01g/kFKAfHgKUx+24Cm5Bw0AqMQzlBnp+r+gy9GdG/AeIEUOvPP6FweJX07n
nKgg049KqXaWjENRL07w6qyj18+Q1OCdgDy5gYdM2+gxK4FK+Qlr7Gjk3CsXyxK7
jzokZw90LnXYHDubIyfrOteV8DaYrkc3RHp4wG5ONUTl+I7Wnv26jvYXmY6A14j+
MlFEp0iVntNB/Ptta8b8s73GeW7OXsCwcHr4IhYEzhufjxx3ez3kOtk9ZU9e3Bhn
F+4S1P1leYKiWD3mEfEkI51bwYWmrcvoj2uk6PtCUCtSgblISdXQskv3OdVPyE3T
EeY+PbMdpdXK1kIVWIaOw7ycq7zGIFg8PlEyMG6sVGQq/b675gpciBickbuo2fH9
job+5N6B8zPSP4fsX3br5CktdpXfF9vngaku5jOOiAedDLusCgq6h/bMl2bk4tdj
zPVvLmTd6LHgADAW42n+aH1DuvGWC/4Ua3gRLbdGQBkNA7gmRDqFH57JIWtTLTV9
N5PBoliLySlKanZf8VSuu/krGsysMBA/FIWYMh3DHWj7w2RJ1h3yPff8DVPMQ5Lk
uLy5D9WCUZlXZdWIxj0CVFxn4G7J/2NBcbct8Qs6h4+57PUgy4bhzlCob5Uog8AN
eQJetPfisIlqwAoHnA9Riw4KE0JCzMMUqA48DiAJlEbq2bCqF6IO38RV/lf876GY
+16DI2s8YBGOy4wNFs/yWQ8Bo60x9bde8fgIqCcUSzvVG+hGO6dn86k479H1qEMI
wzBvLfiWso8SkOxWDqlSocARYp6Oq54jF/jrvLfdeotFyz0Iy+ycLv5Utq91VOP3
aMJrzMBeNVinE6IKAuNIj3pHT16rFZXaWAa/wl/ofy1V7AzFbcC9VIQ+G28Lorob
aMClsaS/iAUpUaUpr4JqzTJH39R6zR6nlJKveM2KW3yzKkmJV4l9c8q5BPGnXkiF
oNkNjtnlG/2LEesq8fXowPlRVXC0guYttcZXo9QJap84TBdcEnABH/lT81+pfVgL
XD+y36gUE38ggPWqOB/TEovwZGbT0z+u8JnfgKlZANC8ardydsfRnGN6camsyrr/
41UbK/7SdsK2TuaQ5W34UJoSo240wa7HR7G/1FnXzCJfIwNYgyYnSCAfrmLH0BLt
Hy2ovEyLk3sn/JaXCRpke0lTvnLhhXl8xSHKb8voI3nniRA2VyHaJK4AstuRK4rY
bUIDn6atmH80dqpEg2xl3QqTGQQPohJGuea/9cykAGx//43VJF6Y7OE2L9H9dLde
tT6UXNeo/wQ0axHMkCZ/nDf/2hdZV1LBPH1o6uCpS1B8c2uzlsom056btRiob2y7
pJprkRUmsq1s8pyg+Crm39qM+Y0ZNbLxyvq8O0eZ5FoVoR1MJl9lxnV+59csnauL
Bw1W0CJHjCSux/grVM5+dDvodlTzDNqrCDFggLDaD9WeaycZeUzcOtbChIlWMHXZ
gQlENA8hL0tZXxQ2b1+foGqWP4n8rAJYlpMyAlmxUf6i1/jOI1KGU2ug8Lxdf8An
z0kTZfVcvGn112riNZVPI8YTy6bNeyH3sMskHY3Nsnw6NhvKzsjzTTfDPNE8HtqD
uY113coIUEtdtKL814GP/0tOtOHMmfT+RQNf9FaZuhTHFZbpf4N8+exvHB6jVU57
1cSCJvCqvD5nQR9qXbeoxUjDKcWg5T1IHEc1QjKY144+GKEjcWelQkWE6pW093Tz
FmK1QglDeskNoVHqCtxDA79nf2YuOt1smRLdLwz1Mo3XgoMUdIdPzO3Z2qD5Jqrs
KAAghfTLraA/HlD+SDpLU7blhdEBVfyOWiXlwaOVD4VK8fZ8WUIhSmpuzO+0+ukg
YUEIHO5rTSos8a0j4cFwWdQxp4cIEzfUApgiJ/wXjjuPwOlYfNdOzAX8v+hrr+ot
x6caDDjAXhpZtNClIqblmJeqw1QUbqtOjMP9NSj90RAQ+yxVYNVFSsQynmyDOfGT
m6TuIPpaPhk2gWJIJrzwsxhWCXrZB6LOrEEY1hYssdYCi1VHZoCOqyKI65o/MMhZ
75OAGlW21Rj4VGuOEA6Rl1W1A1q/dbnSuTf5XaVxsbK8ieMgVmxjB0to+brKF9/z
hWNT1OHAxTyy4V1igzEKVqzpqbz6fbcRvdDgK4HIcepy7ZRrIkw27Khh5CG8d2C2
JaFTiusaadA/vL7OvDqyTidA1MbeF2fpd5UFNerqePpamzZ4q8/EBjbrlsqP4w4g
YnCMu4Zu+Sc3kMa+/7JE6Gt5Q3IG47vkp4VbzV+8MyOHzoa6Jfj+QOE+pi1Bngm2
dc3gNdgscYOGtFffmEb0nW2b3HS5azS+aM6ByNASPNL4UwwerDVDXLbDkgzwVTy5
A+konr35YQCATIybh1CF8uJtGXpiSS+9hrpe7BnALRB0hJypWmDXa2y7ywalGhWx
KZ6bUGc5HHa2cn9QoVrzGRIcJzEWRM95AC4ZDXT+8jKoyMlsPIvfOJIuSg+5KnBq
StZBTv/Wh0XKJ6sEDlHYVW+4gIy2TKXM6M4QxRMVd+BMuycttVYER6wtvgrhom25
y948y4TkXG3sDchrg8Htk2AmMarudvyTa7Fglg5mna0wiahrCldUQ7/LVzF5GEzh
iKdArl1NPmcs64NMmnzTfwNCm4H2ZCHrXRXaJDBrZLEYP/5M4a6sGclpPpL2Kabg
XMufWJSs9EBCmKwEbqoswXKXETSIcRN8wwqSb39CTchd204/m4w/R9AU9RoS6W8A
yMGfuOwOwmZRf0BD2dGdPmplig/Ifle+xwMLLBa7KrqnOizoi+ciLmNuQXYBcpUl
X3wvceIPaW2MxzE7v727z+TyWk/DKGoN3sWARdMJ/KDM92qYx/vax4rJjYrF1nbV
SpUEW6LtzJwQmdM5d2f9quCygF2flC333oax9Nmguxy4CuoilenNgBQJhIe2cW9E
`pragma protect end_protected
