// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:56 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b1u2O9Lxgb+8M3gjJHEj5DJd7pVYSC9bf9PYs4tHgcI+hcmBriFrUbdJERzJivgr
l8edlpC4mHlgsFrDXmoAX3Lc0bzTGWQMkel+Mkm9YKGuMJDSpSllcFn4p53RbQ1p
By5gHOjw9b4dEMuxYEiiVRYepiDpRMzvIfE3H9XLa2A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
EvCn0va0RHGghv7cV8gsRNnYDdH2fa39UMfUc/01b/W5W8fNTpX1QkM40rUfRAVm
+FNizim/q5Iekg/UkCGBpPXhf9xbLmujvSKtyzn75QRJ/AiHpsltlZcB8rpijLsp
miCmnIrmhZ+XpKK6OwvTEjxa1nLN29pzFiMa+fyo2aEP82Cu0lngVgamLbuMOVgV
7lRsfXqNvTfIDdxx7TJmsTvu2zSKwcaTJTavmMM8KzrL2HGuXpMm7zswm+4i6c7T
O5OiyIFp/maudCa1RTr4r3AGpC1tRsadSUgmDLe0S7HEi1KrLjmYreHOcwFO61QJ
eAzI33psyqo0QLMNimaIJ2gHtOCTaDbG2naeJLzmWf2L2zKaPUBVGEeWR1T8BFvg
9hnMP7K7SQ9hceDSdjHpWAwXesCNcRT0vxXIYuoSqnW5vm3xXS+70iZ6z2ILKWQA
9yXpBzOS4WylgusbD4KPzhhiWNaLb6yHIMynnsfiKt4xJwL2vsqauwtcgtsSgAHf
KbjB5A/cOiRLixRDu/mk8QkgZXimv3s6A6HpPLpaT2gp/KN1Dg01WqpgKgO9X1q5
TxQ0ITuFp+cO3qBzchiJE9w4jA4bKkQ5UryUAaOi47YDRlqxmU9Ixr3mkjet2+Pd
2sP2Tl8bx34PYqIpS1mvezlWbQbFdYav4IYsAaIMdyCYNzcJJF6Rn2pxCViORlvX
0l891zyUusH8j0de90kvktwaR25BttmS3NOVY8wzsw27Ntjgh37zfjKVHH07XRnK
8Qqse+yeTgBxXWNYc2HrWAqRW9i7BKwrQM1xQfJC9ZWe/Hkpp6NWxnq4R6bsNUpW
zrHG/1UT7FvAHqOigzCLfsdMVykAt4XIsGa9Ld2sUMF8vEx+MBueXVpMNFfiVzBX
mKr8TVRFF3vlz/Z/KD78n8r7gJRGwTXTzsAfR/83YV6OXjq+/o6ob1c0XRHF1gpj
OrJOrH5fKK5w3oGQWLTgSqJkADoi541mS4kb5L+s4SSgu3X6mw0a4nz7YGGpSKF0
umRH/pdvkjTlI7AFL8CNjdZ8oMitcpdB5IN31eoDwS1p/TlsYhoW0tdnktscjdbV
cwg8kzbG0XYSYLBidNugt2F6r2o9S65VTpVPI2GpUj69VUD17F6grkOYCcFokDjI
8w18TvZ7wJzYP+fSpg4KIHrJarqvqmOFdBEFHHM7czgHcr2zBEn+o+mgn+zhBXK5
ecyFdOO7vyBqITaGpf0o6qa8lwH+I/Ifnc+XOTXqIIw3eCc++vyEQH0QkRDBvXRx
ih6z0iXrKunMnCNaRFPS+xpQ3vMk5RXM8OJzccGi8gJmtawvV93drIHXeBI0KeRH
J8ASZ7RBapxsQLA/eLpQvAl2Ep+EoBCQM01KS4rlRnMbLGu0inrwFWTlLjN9Bze7
XMthIyg+uBUGCD8B3E4g01k70O2rTT1KB1T8g5ukOhdAMvMhFcNn4nm55Sbez2HF
zvbIzZhTRUYx50qhR9dmu4rSh0X5X3Mkp41UboU1IIrUdKjT0dumfsaw0/aexMF3
QonBoCukcFXdG0yV9iPdCEvskbX5J93ewnCC2WfvXluzMUDETOdgGelvJCpTS7Zo
dsjH59A/3bfOPpRtWXYw4/Ub98j8GvjCcBrPk38heLV/z5JTX84WgiP1LTGyjYvj
V7s3AKOBxkJHQXLVWUaunx9J/uZQH5bx22Xp98rVJwx2ct5r6EyLRRcxANuoa6BH
K5pUAQUJSpbWHyOO3YPoane/VCGjCBk3j3/mvyXquf7ICGgbNH1LoSJY842p25S8
upnl58OhRIYARvzqB4eS1h8Z2cdJ3JTd4xhovRqQ/U98gVrmWG7iHZ3m8Sv6NaAn
1QCSZOvRU8a9SOCWA+81Kx3reKE/mbjF+K95z9sE2DMAV+g3QBcRmqxGnhWS6Ktr
oxttNQT6FqACWuFeJ39rjtjofLG/GtLzWykNrl2ugJ7rka9vRSWcOGXt2ZpDxCrR
INLcHFAgaqJwQ4YQrjvs6c4176znj4R/91mZ92jalqz+23tz5ltke/WJo1Df8gOy
LS1bMhnqegzyMp8q7kMiolLxgh3k6sr8gQw46xabVLp5VuVA9pkP8nk4hHVysybA
ObdXpPgB5ZGGYmzBtBR7+0gNbgNT4hf/NVJuPepaYgmvf9pKVVHQEtW6OfZLR85L
gv1+E6Fi1EzkxR9/faKfuTG3+WFB+MZKoaiM9YGFox4yDiK4mW1UOT74XcxJ36aO
UQZ7Y3AIFB2wD1DophxJyKZKPyuJlw/OqKhkE+YyjIBGi9YsgsfCdZVt2UJzmIA1
tmdEbnR2+pyWS4NLVv0uenJ8k+aDEFBtIHEqQ1YhlvCHBU+1Rfnnz6MKF7LGik+S
O6WGdDu1Mnu6c4XMwSVtGe9qgE3rezVQkVsV8K/XDLmXUEXA6sVztiUiBqvxwyAW
6OPuy19rFi9owsfM7qyXkGOsA2CZGK1YdTgTMZEVrtPfh7Iy3nalm+gNmvlqszXI
Ujuv1a5U11Udi6rGeSm8HzO/GxjT/KUn694agXlMuk/Z3Y56IIJ+9KfDynSY6HuR
DFNary2ug2FPIzvJzSAhtYABEizbXP9NXg7o1O/J0CDmUCRiMfpwIyXTyZWBRDX5
dU2AaN70aoKB1anxeOMChbrbWB3BSlg5rXuTVkMAYK99L8gwZmZYumT9JmyAl1/G
aoRKUkR8TQahDUwj7hHRKKENNBQr57TFgYi0XXdS8sMXIUiLnVMzwz8j3MRm1iVH
M8KpjVCyxBDn9YqahyzIUQ0EHoIc4zPA4kv7VAB/YwT+bNfuNKg8oT7B3WC5SBFw
ZHYUlQKoFQQO/pPglm2f4eahygbJr9qnL72rf44JCvqhwSsYcmt3I6N5sReS3x2v
lLW4loIGrym5lalUM6SW26RC6pKGhp6c7QaBfNhYtybyopSQponqCQo5uw81QoIY
a6AImEFu0JShSHhF/hXtTmOYcwELLGIBA5YK8WzLydcD5O2vG8FlfFIbFGFanDWE
Wdx3HMz8iulQ5QLA0QUJ5nNrUuUPftYegexCxIKx7PmaL0+4opbONamc3nzwVDdw
8YzsWGgMqNwDidWSBRXcbklTKU2Js2VIr1l9vzyoR767XkgZbRXXq/uTtDUGIX2z
L35B321yFd8xCSVN/ue3R1dfVWlE6WgyIHvMGhvv/Pg8i3gya6/QfUXREupON32h
qEs2m4FiDzlFAenDe2nT3A/RVrYV/EShL4e4BkpAe8Z0BgBL+tKgTWgXO7CvzCCV
goG8rn5IVPrf3GS6xd3v4mPCu86cRjjr8s8V0mh0aiZ3H1uCGy5//LOR2lTnuiXO
rZdAIarBp1CkV2btAHzDQo7xCPhJZUz+mGqxmAIl/3gSMpExXVKpc5pqtecJ5jrw
eQFsbcaIHRDUe9cDEZJc38gB9/FqT28f5DNu15Y3QC3FWNFeIpM/BWGtcOuZei1V
v9WzJpD0wgk6R0iqy0UTh0HYEDjpxfskSwzOLYAzp8mqVJaChOa5PMx/AQagAC0G
/8giKwlJ/kkslXDSfRtRLsWOk+1E08WCJlYCuUGoc+SsbRiB2h60Iqj5M9LN6tTN
0ZXWIFpkHwEnLGdtQTvu6RAKFewt9tXU794zzYL7Efm+fETz8VR38zOgwYMOxfkL
TV8Rojip7uHdColKQvWlapqTTu5cNZ7lSsU+qpo0/LmRUzOSMqAf1KzaOXivRgIl
8uqHa6x3m1djFvWLDW7Xveo89e3iWsDXG2y3Spod/9+I6slxmf+iYSS/eYPE0vQ2
eTqy7P5JAw7BzqOQ5LjVXh8P4/1Lg/pANZpL7dWDWYWQMdioIv3C4+eyi+hBE5dv
0SBl/zd0HBHvm0KZUQ4Kx3357qZpzBMhsTUGEwR5HXkZMCFm/ixPQ0Z8zTb82tW9
kYamv5wX1elrpltkLGvjPFY+nXM/cecEsoRxIm2IT1FAVCQzbfTuk6WiX2fH+AWV
t78iupI/hGJ9ifqvg5qDeBp0A1tq4K8tf0d2LZbhNhaFO1mNMs19OWbcw0eL2fyZ
5EtuM4ipzVJYzRrPR/5FS/Z6LXfuFztSGFsAoJ948coaoWdyS6NdgJv2UMDwP5uY
CuJg3dZVuhWc5thXlLhqnHFCiQdrSZCqr9HCl+bXj6BMs4sVNO985TU8Gqrso3C5
kBBQBIuVcs9Mj8ZPJBX9Bym1+EP5MIMCdgGpT5wC+gEIjw7ZxW1c9DK5yPG8HxFF
qPoYQXNq3t0YF4E00BqU7rJlF/hd8OyfNKUj6+1YpWB27hNj0Pvod31UlnAND51I
fKxIKCZODJdgP4aO27CymhxvZwMcgHm/nzAJLAaDKW0PkppTWQ4GctRkwsTtzSz8
ywlr8btYOw+ebE+80zNhZDG0Vd7hlh6HR9LdrOnO37w+QMDWyh/agKqlG2eI4j7z
l2XQ2HYcbvO5J8qez/vhX9q26QDwFdbt7Eqbo3/V69KJS51Co0/ntkktPAeEg4GG
l4c2rPdjQcwOjHF6xGMT2fraVh6+vIgn9B2GfOJG1c/e13KnQ4ubriGSMP9CwIBK
lwG0YZgv7zTTq8X9LI3mgsfqt6uSqKcljrL0+dI3R/LPBBrOQ83FduDzf9dojpnI
GFDD3zppevIKnp9FYtS+oN+P9zqFvTZNVqZX7Rb/aRSY4p1SfivKeR7jsrV4W2jV
GgirYCUB1A7MZkePGNVZaDgYyahJGyim98LB0ek6CDkVUpigo89qmH5jqVfROW0r
dy4bOpV15waCjAIfzO96fgpjT4RCX4jPSR0MU+xulr6VoFr/dEI0TBxNg/WOAYBU
lh7r9m2A8X/1aaQ4ThBXUgXyGyYkKxRt6yZ0a5IBDqr9I3/EvadyMF9I+G5SF7pP
NJ66q55psLIhCtFVwISpq0NeqqBtbPedjzoYS6GJ47BsUxUNyqeZBoxBYioF6lmR
lrxHwwCQjBoIPmCTK2KbZ+0tFNHkcpuXeCHxqPuqxEMDmVBqWwIOHb8IsgrlRzsb
JuyJhhrWpV5mXHv3QLMSxuSLr4ZJQFbepn5j2avmNExD5+ZPMZRA4lJuoelEfXaN
6Tsqzm2sxR1UBHlBCMTbD2z5GgH/ZfzTUJ5tvcd2kKdwg1wgEny+FpKNrKT8Z5kt
2pDYjnS3WtOQB9qhtnQUAOOX+gB3w/CLGoW/ywDM/aJAdbOlsgg3D1gPaycHF1la
ZWSHzN2KWRrcRG47peP8x7uqA10dFtBd7zf5rRpz2fMC/Tvq6j7YVZxk0DUTG9YJ
m0TA+QUzs1KhLU77Zb4eMjPklfhbrixo6BakZjABwfMOp1gpEzoQu5wUV52dcBE2
MDYWdBoKhvi3L0UJ+vN2yQu/deezD8uEshVv/lixSq6RwsvDWN4bFgabxvr+OARd
QLx5/2RGmrZ4e/2uxh1r0QYpj6T+cxL7PGmkZc9f+do0qyvTyl6/vYTy7GJrlOzY
LaVLOm+Li3e5v07oydQ2bDqb7Y1SDv+RVOddlH2SBReS3mP2BhzLSzllaMtsqmC9
97EYEwF/qERiU9lNQ5BXBUi0Goda5emME0A88xwjiwRt/HtuzXeRSSHZ27Av45IY
XjYLzCl1ZtoGg/FScZULhC3PEJtxJ6AFoSooSmCoCpn4dd2vts8rP+MjjcwEabqS
PF11F4zyuns6bfqv+kwbuHNV3zs5S+OK0G4YOc9wbxlKkrfhTVZ5Uzhag8eQXcCo
cb+nyzQ685Jk124iuH1ncNhYixP1CM76q10jRkIGJr9Qe2RVNJR86L3UPIJVHhFB
1KqZ0B4S3ciZKMbrymMqYGdJ8jZ5YRshVakFmeBFAnRrc0FbI/d5psesSYE5/p6J
TYEO1erwStteaDpVlNIMsVISBYBEBP12W2O4RZlDmv+QkUrUEVNGr3QnbnPwJcRa
vQUpn4KflHcxKwtGI6nmkK5+TbE7ad8qggIl5cW2BvzDT/0zIBwwnc7VUdNSx4Is
NsvQe+JpFYoeV/8mchjpKMiNVpbWjSx9OgOAQXIVr8nm2EbCelx+JXZwsQoFo3hw
GmhZ0M5sV7QQlpdDwHTE8hLRZT9IlbIfp52gbjL3MyXDS0qSFuumC2Pc0vqNdaSl
S1zc6XxLTc3XPkeDYfT+TvVyf39jXnYs0F6oWX9ahAsE1JeeidYY9Ty2J7uYZvT6
RB5goSpEn8b9oDRweLwgY9MZV11C/RH+hmYlx+asnyOlPPrby4zUa3wzoIvrgCEi
NoDMxr/jHsrXFVfzOyORK2KilLa+CuXq9MQrjkemfBhJb7tMHCVyVcKmGIcxitrP
iwaIy6KoDpEMiyrosO/3Zz95tU7RMN8BXVkI0EPky27zloB0dEOZDLhatZnJskPv
kS/D7lyJpWP2YOXUbTcJYowIcMfid7XJtUKZOhe7Ynn81777pu09UomMw6wjwt6m
Tr1jKh2W2fIG3ns5Y3+zmnnI1G5Ng/xqNyzUJ+vORYwwTdGnP8zxZ7fofOXurlLk
CthUxrch14U7xt3RXuoNf/IOGbKukdgZzD+E4w+xjNVWql/Ts2xvqtB01o29cMCK
lqoAkBLQBqU6YLjxsdbW/MTKGQ5tWIDemgrKyn6bNomQHE2hXmkk8JxjUZWc3aLL
+PiIA253Epk520r7WhoKxBrCng+DzzTO96Jx1oiO8vloaMos+dys0ELL9enefKbc
ref1DM4P+aQOz33ZoB2iPP5ZCc5hrmy4hYW0HYy7+oFQE7Je3xLUNY/Sh6gDO525
bWarAU7Lrw77PkYrmHMwOmUnGaHiGdxkuttpWPhh8s4c0Fq5dKeKXV20/vuiXmHb
atHuCiixtZD7OLQGitFD0HXFZWYTn/VsEZcxpAugsYabcLibkpFVL5QyPaWAY6xc
g8ygXfycTnyRCbnrcgEIFvrG21E82y811vwTStLdKnLXdh3d2dXDckl92oa5hRre
MbQOgJsEz6zmJpQcAYX72CFqJpFsKx7SmHayl9du3yqS44DB3fchtEbPTY+HX63t
mqfjp7mOh3C43E6jUQY/4BWG07GbrFaEi0TPv4oGy5GB9Vop5zAZe7nU8ASOja3q
0mKKn6196/vK2yRyijaEPkB683gJt/SHaWXlM1fcHc8WCvDAnWifCGXfAG0Fz5tO
AHmPDMaPmetihDVuw0d03BxVnCjFH2gn2Mg5zsOoyu5ih/lRocHLfqxeMHnE3FOw
kgNkU3IDrUhO8wYYJHv18+sct9qp65PV24tF/LP43bcogf1GevAihby1kF/GyjyJ
+Kl1LyDsnTr0W+l1Kza5zmRRJTgD1uvSUx4jXAofFZOAQc4Uc2en2NkJEaYFW6i0
Jbw9572DqBCxlkDFzJOV97vt3BsCJAKjIEElujU1EgMIJZDUbwhEDDKas0P+gJEo
bjPW2pnPJc8+oqrd3BFndGv58aTza5TGxVWxZr6A9ppSbZz/hZ946pLvVkKL4Aez
62wfgRwKpiny1/7cy8Fe7CEw6EnRB2R9xq1T76mUVo/oUl1iiZO97aQ4uX7iI33a
ACCUAdBwiGEae4PZBGk1ImgfGv9LrjwupG8xA+tuG1WBs098RHF2FLps8x21TeBi
`pragma protect end_protected
