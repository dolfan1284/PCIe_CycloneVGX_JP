// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:58 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZObptnc68FMJW42Ono7HB33F4+svp5KpYB8K6ZQCjbm9U8WBr590bFd/Xf+ryxqS
Zhs0jRrs7fv+u7M1txlgDdg84XVx2Pb2kmJSTPdpiFLVRSb/lyBVeGlg5xJ93RhZ
DxvoIq31ZoEynA3V50KqowbIvWwx9WwOQ4s8wz+B2GQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3312)
XWMq3NycwfffGUtf7PMpvS9TnWIlc1BpkitdrK9scAY3HkS+c5yZuyUj1JUjBRWE
UpzfoNoSCWECLjZBcvlowdMkFCPiG/oc3NYeJlPoE6JGCT9zLb0+YDOaL1Q7569d
F86knKKtFlWhhAPjKBienGp2cYETcwltZMXYzd+3y5wDdFfX+TMOaBT4QJvO8KUM
qHO/nEcpIH45+sSRRr6UVlN9TUK0MD99SeWRHV1eqE5e+Ry4BdmzP+M7JNbbhZuB
nZnbqGmnsLv1j68Y4aFb8ZJadoy4IbieCtuMswOILbsYH9lqeenxB51MSYNnZovn
zFDPr88+JpMcW/QnwZg8Jv510stAU7o1Rkac9x2oQig7Dczx4DXpjYZlqQL7grsN
HV32nn4o7GEdETD/2dqypV0RQJ7GKuMfe7djySsbHXnUaaWPQwjZOUeZHq3c7+l/
ThxxZINjYf07QQqCc6yq5XLy/o/Xs97ToFAdG0f+bZIWcb+crymCnnRuybYaEeFB
R3X2GY4Xw7F0b/dvUWBl0hQkqYzP9TJd2plRBzQP0PfgB7sPVzYcoswurtVy6pgV
Pfb78pU0gN4+ezRvJI1o9BRH3we3OJqf5mH5jhyHm5TKGihHBMvtqfM/KVjrpbh4
bKJzVvzCL0iOtWQbgapAvyaXWDenq4dWrk+K8ULrdCNPAn5ddRuh3kMpk3XOw8E2
pKy9wjriYXEk0TqofvNtBMYiTsqVgvL6EviWwVFexOTB0gMdMR+WCNHTPA4Kt89v
wE98VX4Cm2VrwPE7p6bjJ5FUIyj5XWZZBp2GgtxEMs44PW5ywnHXN8SE5xQDvTXB
zpbJ16HRPjwxJodhrNIll8O9jSTZSxypI+FB+jeFAmHadR70HqViCcYEfzhI7bud
EOpPybT+6pot/yCMIPeYSi78YOpWH6XF6Uq9bej3P3xKsUD47MsNj33cuX7AfL7a
tqwxTBuRD1wZKgsvXQkR5DSh/aBKtZIzcyxY53kscKm1HN3VSfb3AVLR39Du/H4e
6QpuMghS6DBAB127DsD3kUHfbspX61EoeEOP65L1gr0mbPqvoLBBAOTQM3kqcUzo
+9imsqp8QDXkWDkGHqBLs/Ij3cST/UmHxMiPvq0t4xiMD65EeSyYY0AZYoH4qQaj
SUG6NUoPPo9UpdxtpX4DWldGvM2Yjntm3V2N4/TtJ4313NRzinrc5zYMStZW6CL5
HD6KAp0/6T3wFYWxB7/yK9g2LWnf0J8fejp4iNFVPeo06mnJGnTjeAoFZJplZiS0
UbXfrgygEzoNRxi1HsbMicWGg1PT9pnVnyn0T80BVcOGS5K7TcnakQQZnW9q2Pzp
rlHru/eNekBqY38laj+Tjobc5wzMGpyU9H0tRotqjJ9EVnq7GHJ0OwQwAe05Qjgi
cgsDHqbUQtx56ch8BQNu/LM9hfNAAoUakRNMXZeuPt5h4Q1yKEadjJgtCxAHJgOb
s4jQtXWvuxdHm/VZTj5muhNFUiZHL5ZG/CFl39JPwVoIvNQu4h5UK5c3QMD8iP5k
w2M0b8KOVSSra8qxWsgWYHApcGWabZ9vEWxrGC3BJk4VTrRR2upG0o3bezuki1mc
SbGLuybR2Xyiuodi9VyScr+XbY4sRE5hlS2XQe2pE5qBr/tE35B5gcF3L2h26Elm
C0bg+aqfupkVMHlJZeTAT03TjcvaaiVnWEaV8x87NA5f8vdYiaLenuvQFhlmt45H
R5tTZAT7RJKjU8s+pmsnEux+XTpa+E7nCXN1e8Q2ak1NktxKXSkbeN2xtpnHW8sW
Bj3QH0VpTQW0o70hNLN0M7nQEW70OjTZa5SDNprAqDWP+AGGkJC/BH9+bKZRSDYN
rWEZ0LcFgCmQMWHD5d9l137JMpvu3CN7ISaR3Eb8+U00NYxvIRmGGtlxby1SZWKG
Cc+Rs8ScF8aWwjv+niXTMOE39h7oS5mPosX6vcFKADM+pTe6Eb1iTFaMHUfhXGBf
WMMegjj+VD01arFZR8ajJZBEQlbaeGmDCJ0LDIrOHqgXkkXDL2RWPN5+cAvZ6Mvy
TBm/6dKW/8vsAcGhcEeLvJLzgsl5u+Tl45Pj0NFOdOOQHVWaGqeJNWB5ar8WEvZ5
zIllfebQaHddiczpNXMGk5JtA2Xv6qb6cE+Gq+E2VvvYVUPdujVGrH3e+INTL7J3
Gu8RVhjODMxfmTEZZbn6xY6n/AlUSrLqw2vGH3qdQgoNpqOJiFqYPqb5eleJq9YA
m5Y6TKmELBFO5Gd81yPiha9RRa4VVGr8lWIZ7ewcLc70pLTB+p29h4ov8nIrkiZp
hP7Y2HuYSXLkCFWzq/wzzDHeNE2SRwsGu+i7VSeL7SlOA/LNT8qQlQgDs6fugQB6
nHjx0Jbojq3rI1oz+2ttxCnxM8pRQKc3WWw0vHD0wRXJ49HxCt+hB9biuKQJGm2/
4xajOyFLEEbwnwrB6cU2CThzojwe9wFUq5p1B0e/O74iJqJbH/gvbnkhtclF+BSc
q5mFQqG4OvgorAMewcbGhOa7u137mcWWhgAgsdYKJJECtI4OoLz6joNRIeGJSpCw
/rFBJDpMCy0webXr3UuXxhqkFhspAytr62pGDDBQHWEYtp1XNr20YMId9ATIMrG+
VF/vDiF6aqxoixyd+t6wx+B0wOLp9R9Pi5hZEWIlAzvRVfjZmRW55wUL9C67CUaM
RsGEhbJ7NP0jJ5PR6c8iVqOPbbDfVZH0K2iCTTx/6rZz3J3zZAg1lkSirSchHfXk
brW6PighS3cnFFozDVXl+tJXMJlS1fra+V69oP9WslVQp8FevmskVa0e6nixA2z0
5wQj8X0gkCAdDF6Naad2gU+s7JTyatuZk/9UbK9ZqFdYdBbyUElr3bDiv5zUGTEy
AXqxRrOFyNkAE4G+40qCzbW+y+ASJubPnNBUs/UPdAbUVXajfRUVed1VxWRWH90f
4zpdHt7yIZtazjl+NKzT/elXGkNeRn0N76R3cPM7dmQiTQZu2mRAndeyRWRMhk9I
j++AFoPkMnvsNCatShHCU4f9OtlJiJg1mZO5/iVED2GnRZRuzysrsCramU7X23hj
fUVTQFoPZ61+0hiGeyug7h8FRgpn1Z1oc0XrZgHCpC/RgPYD2DGLl4GOo3llbiSp
0cPccriIyTFRIUSQ74bUizkZTMEEd3x6vTfvWURR3ybDjnQGLzPKtJeXgLH4TCgB
ktGsspUNzKZ+AxGRV7bMpPjrn1npx69ZLlwZeggeC8K9szyksHxHSTn4Y7Ub46Z1
zjIt5MBgmUsYaW2iWARZGFmBrqvtIiWwXPC6F5Uon2W5+HEon/HBmu5PtV3oGu2z
IV8nCgxxvpqCRIZOMLBhfKg3nofQcwe/WaMWuXc+5OTn8+Zr69unKNyuilCMoKTk
n+7S/rIuBUwOXN2geBXNIiWYtK1vYeAqfvqeP2zKM3o1Ede+di9K0nmHk8OL0gMw
DXPjRW+eMHlS0/3+Yahu1iyVVvCwhyi8SaQ1pVl6mCOruQaRkiLOvuaRQPt+uFk4
cZZ26KXfQU2o1yMK5/yQ8Hr21IizZnAcdq5/RBDm2hju3IgQfk57iW8mPaeeMiA6
0kqm6+aUaXobBEt4pdSoo+LdE20YPULh6vbD8nP1yTYDnxzEo8C5IUH6FL2I5bDs
rSS7uotgHhLDyFbX2QrP7HomC5k8g6ar+ih6V2NgRpF4gZ3XR4dO0o/QjdAy0Mjk
N4ysHT8Wv59b/KHFU0bQoElDVlxh581R4R8/1oP2bxxSEPzvmp64mvK8KBgW2AnN
ix7DT+m7qr7zFKBJL4+XB2RCSzBXH+jJCBPvtJ5FuVjz0vLJ68Ax8SjOpVRqDQjV
N5bpuiZWpEOrswUC2V7wYpk/FtttWsp6G8RS1xD+/nevDQ4uhcz81qvw5Tvb3/w1
fE/gxdwdOnOsAUQWY8V+yJ6N0mJZ+U/3FRP2Au7V5btjKXVtXaEwIGwv1acn/QE/
62uxRbZRjxNkvDm3Qqjx/Iw8vKxjtyZBEav9zIYmCC/C1ze3YwiRDo4zkei5DHMI
KI/Uj86cfZC6wM8ES35vMPkt8JCll+lqp5cE3YwX7WQSCR2EkmFp+HML8KsDqA0h
BEdLYsFFjmm5iofCJZXtD418GoXbPSAUEJrlk5Ip9+MmzbCuSDn6DvTLME82P1Bq
eCRb+lDKSUnyuaXm/kyJXMtOHzarrgocBPcxe2b036QyoEyzpdh7uf702/9yHwJu
sqCkPcp+uxl6sYg4PJcoHkTvdGGYmcGoTOHkuF2ElacjN3Lc6NTnQtp6RNe2kL8x
kbRYH8UZdhCXtLBJdnR+qCwxE47Nm8Dsve8/NuSLUSg8nu5AfMzuNHbe0l2K0i3r
N8vOi/mfbssQaGnFkduo8V6HZDc/ySPvLyGLI0jthgRln1oOVN1Ivs1l43Woiiw3
`pragma protect end_protected
