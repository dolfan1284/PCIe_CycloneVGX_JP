// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:05 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BGVxuoqlWdgJPElmE0HE8MNNGqZ2vGmjm2QqxJdFkw3KWKTcD9VbWxegQfUGpuha
QJGgKp/8e3dG2XPmHoKYECEt8SGQmY+zQxpmG6m+ZMQmpjBRaPja128WFFveVu29
8PC8pFYONyrIIv2ZyFUHUsV9zW5/4PfzxqrfNPswwi0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16320)
yY34vWt7bKHa6NdhUzvPrGIzHsBBT98t9uwOvsTT0Ng2M5EruLQM6GKaFUuzzfyk
7fEqjbA9DTAaGgLwnrvn3FzPE9EoYYUDEAUYfB+Y8Uyrd/BRlHLBT3giq1pYyA9K
nG46hIDcTRs8Iwb+v2Ibj1qzT5LkM/VyuZFgA/u22xFeQ+cx/j1WG8aV0gFcwAn+
hBM8eEZ6HSzjdRRWXTrw9Xt+kOU6EdjJ6rI+b6Y0+Kz/Y3gOSVSq4tRttODJcOAI
IMD9F+AtnuQJrVNjsu1Zl9RH8AIyw2cpXKbVRe/0Wqe2qenuSwiuysryF36a7ceV
HcgBY5yT5CwAsSudyLMN52s9z+5O0jCuEGr7DMB+zRlN0FipBGp3nRJjZ62E9Hy3
FrKdSFfIq03g0OJ/+/szNiIuhM4aqRJo6PFNX2LoPftPD0wm4nSYfHLpEMtFIenU
62oyKYuYmNyIk420i5K6O2TAFII2blxN+s9PxH6YVacTZpJ44am9gtW5cgWAQrj1
68cPdZ3w+ppCHuy/KkFenwyKET4Htn9de4ei0VDvvSKKIjV/VuaZHiS6lS+jRhqg
CHVBAUwo+HbSXgBRfBCmv18BkulngRzBQ3GWQ0aO4vGt9eZQ6JC3A/CEKGfvznvA
8Eoy1853fL+NBEtk7zJd2ovUx0zxIi3k5r/glT1eWSEdkDa6zBfNiv1lMRJaEUTT
DhEdWbvysM5QknJo3BqqKIGtAN0lqwVWJAVzuB0sinPYu3v9nDl/toljFbJ5Bqai
SZqgshdDXMSRt8s60UEcEr1H+Wc91TP+u9CH2B2uGcyVDG1rZ9Eh6x87du07Gu8y
WuRI4rbz3XsZCTQ5OSj93f8sBfe+rbXbyaaLdVZhaDjd5HoYpNOXbNmTgavG/HAe
lZBlf9UXZpIbEDNL+H4hfMAnJM2gTxkahWRxNj7Cyu5EdctysRjdmp9PRn59Axri
yuiC5Z4ljYBvCjXzZmqBwT1mtWzIfQKH/2hFVQEr2PQaiIM5bI+KPJxNe3VurXzr
KsHmTETdgQXgsyjf4DU23/S5wYV93LcVLBXAGgkVqJ4CrXhfClGC5D0qelq/2ydm
WBSm1MhbELCVe8LUURKDc/RTs7Gtc/5r38wYwTOOujIF4NyschQFMTvsFHAzJWvK
d6wl0VzSsyLe9Wg74/LlZupRCPKthwx1T1GkTH/7gzknDSf+ZS5n7Qp5j2K+NqLm
MupNl9dm1kacwW2F3WuxV4bxpemprvTV2qy7jh3I3DuGzM98wwB4hL5qrpXC4tuX
BGMGoBG3xN+9Y7XUL9jesSn6PwBnM/1sXAoBI4RO5LHOdVdSGbo6YMqKpjvguOxy
ZNa6RjyzWR+91tj6+sOG97g5LlGJAsCvDQ+WzqdL9nBkWQLVYkJ6qUZazY7JseIx
KWxwHT5WKkWTHm+9T/CnOuWt4vl4qQRrAQMR2oG/hgSNkupJ3nxSuGNZNgIWJq6N
yP1LVis0rtO8EFCe2akqsWeElUJXAoxsl4H6aRdlWuZWsJ6XHp838iP5GtmiAddE
+2kOnTv/rYvJW8mRR3VFcO9lA7EPnJvdiGMTDH9mpo1Y+BwL7vVsBGGHEqqBJp7z
K26sUzve/BXbhvzrCJi96d72Pvhzjhz/95LfxuhCEJ2GJhqdMlPSvRGZHRk4nwvh
qwRG82ybp0kqB4+6c5JsDI/dvmS+mfL9e2VWMixfeCGU46dqyKt5mrV1yPC8wcEs
nqL8DzIcz70AdfPnBw6JioxGDdCMQ+pLNN6e5L/h0Pm4fdMV7gZhtI070fOZkOnT
dnkIwX7gZpb38TqqTA6i1MawN4wud/iur5ou2oYusEiRq8uzD7FQv1gZazA2WNkg
H2R8BIF1G/B+3zA3QLcDeMnQWWewDsQaLQLIs6hI1ibga9+yDJ528fzfBtj8qwFD
f1R70wvpjzNCJsmVVn9VjB4zQBVYhbbEUpjqENMlfJZKPuMF/jYWGqJeYPvQEST0
Divk/8irXfVcAxMDkyTR/QeXzIU6wTcC3jHoGfClqJCMwJBNWTODLdSmZaw5EpRA
D0YfBKlo7f8t/SLBqAT0CnOB4DHHnKQiHEGqcKoCRmT+YhfIXJiaTc0xPbmDGLzw
jzs1P/g5xw9nmVg22t+MVwyUQp35661XBUSfH9wMD1S0p1aonrb/KOIMXXzCcGIi
Mw9nRmALzhKQjyczo+r3JxVYTFvJTsfBLsG+GGOqIUbBgNfzU4AxnyNsYMNeLVM+
zwn8o37Cmx64ajN17Jgg1n9RoQt5P6NZ18idktnm1BC4Z72+f2LvuqqTG51l/JpQ
zAHovIy3WJ88KF0K7lhO/w8A0P39jBuM6dzi5Lk67PfEdUDZlx9+XGiIZTTgb8UB
o6CQSsnnPMpcvafkL8DiVx9WDdbfukmDmO5D2e1fxhlvw+WQcrvNJrlypIA7obv5
jnuc82JyzEuyEBh57UZQGTFrVcYbp/cWbC2/UUeIFd+ITulgZjSBil4grsErcgDo
UVugj3m2IXPg/QKgbDc4bv+zGyWjH31OVZsud4Nqjd+y/I5damLSDSSO42N5qaLH
SnEZz0hTXFDlrK/lO3whq9YliVDHOABgM514ITDExPH9+Z/W7bhxwrSLpjHDxdE9
kPygNb4RIkL/nRqmhKD18Y27GT0FRouHQydb8E2GTTe5QfqKJh+7mJyPESYxUb15
KSaHbAYAtfduetDHsdt1RpQ/9g2qi4Rpo2MuCk1QaOs7KTZcKNzJ/HLxbMaWd9/C
vwUwVg9yiVvvEoFcqLXSsqAQ39FLNB9LYywRrdwLo6cFgpvPRiuNEjKDyqxh5/AC
+4jasMrbbdvgEDYAWTcUKF7J+Y6nHeupOYzeGMbaRkGBTnqovMUhyiGA4N7oR7nX
Z8EcRFBplTuecHmTS79s6rz0z39yYvfFbnbugAVW8Pnuzcwnj8oJyGEgmc6PGBga
A13lY8AAQjp5dkn0TUWnlnjTcSSQxyDS7hWPoIv8DxIiGCTk2fJJf6Mg3jE0xBfR
3926Ih09oOKXT1q2+gB262zWsAAWvXhD2Wv95Aw2mbLja3nq3puItxYB5Q64srJ8
FvbKchAiOZj0EFERe5YUP1FEWA16hYxyJCARsOlT1Zsg/M3sdkunGURz7D7SLIbb
Msd2jHK1y6myNo0pyysjzOKuKALkSaBmpkrBzk7kleNa5Lun6KbT6+ZTO4QbBOdr
6W7/ia5h4VMdJxPhvjmgTSL49dWp3n5sQRHL+9cIvmrsOFJrA2HO8OZFCREr481b
uXF6/OMwPyC+9j/fqOvGd6e+gTW9mYLb5V2FpB0cJqIvYwZulnRCJqxqtK/tXiwh
CUcMOZ9BjNGXzRC2sRZDm/98OtY3SeTSRRAl4DHrMaYhJeWaayLObpOPDAqpILUu
BDcjWJAghkUN7KinRBEz5K1Ojxf+lG6ffwYdF1YlECOg4RKE2aZ02FyKhvVvC3w/
k81zBcgXSWaMsxfwrWP2CGHo1FDm87lsZ2z+yLs0ojok+bPSFijPlCdXt9GTexo+
WJ9Pu68fdnIiQfylwN/jyLAblD9SyrgHboLX+PFiraa/ZruJvlDVWKmHmIFwXpej
5hpQ3sVadxyRnCgkY85QGe5RJIM+hN1ui51YOpW9hMOHaYtpwtAkKrjAjiUGcT1f
JE+xXE9MSU807X+QIYNEWO2nZmEoNYxM8EBLocam6mA+hv6EgXaWNCq1wxK/nVih
GzRjpgnMtEmmUoXWykWQacMdqNR7c3J6w2HMp2vSWj7I5lbn73+vrLeTqSCcpL4I
0ISq0jYYN7aR60WmbOk2qzs4PohgsE9e5PbStkMrHBW/MZ2yPlzhypBsocIhFX4p
a5duPc3uoxat8tbumoa4cNWaMr6sOPTqxTFWO9PW5LNqUrCi2yQ418xFearLrwK9
mkTnEs8IDmEYsgAcrceeRoXq226leTMCjVTVN+1B8cZNDyL98/FvRttrzBy1ACdD
Q1Yv7dU/fmSAflU+VjPLhziuiddPGJG4CvvrcA94qg5kG04ssVm1N5Q98r/NZ08W
UB1VoRdSWXZmSrT2s8Jr0WGyLavQBIqDkVgkLmbIXdY0uPo7rqO5IVYQinYs27UG
mQ0rsmVefb+JRPyZkg2C5p94U2cdbe77+fDxkHhTykZ9WPA82/g4XoBjzMKI8gjx
7mdbjjFqaFKYzaUiEe7EkEi5h63dcnL1ahsc7KD9HKPwpyYyrgk7Fw4PDEYz6poy
l3EGjx84bp1B+uzeXT/LFKRvO41YOTbcfTtesnIZmeLg1Q7qGiInpNaiSxSuOi6A
U+2OjJFSG4yYH1AIhi4Py9xQEXUELLuzz3HN8Utari0xf/b+h9N3T29P4/3Xm5BL
JRi8L4CZYvBYnpYb9C47V+yptRbmqFg3qAFcii6qrDGJlkTQlFKjp/TMqyiEAxrt
q2cOAAFKkLR/2qgMK7V/TjE3g4Mbxkzjl7xYoNHT2YZWIloU/60ZL4QpVKtKaJhz
akmHdG7Fmu5TQ9KzgViEHP9I+EZ8OIz6rFGOMQzGzCcCz2KmXuf5mTf00LwXgKbx
8pMKMiaSMzRMmxGg1Q3nPbrwwJaSsi3fb87kP55tthsbgvqbdBzG9+eRZ31Iq0DX
CAGWqrFx9J/+S2L6TwVToESruv85wqnjtGBDzoktRED9inzYkF+AWVEgzSi2EUaw
EkCEZ4W6BcvKqpsugbMiral9EgxrlrKyLrK+iZoh+sLacol6y9K3Vg+BE1fw0StU
3hH96+/l/PIB3j/62wUrZ1+CSgAkVia9VWY0CCOLjiLlfR4pbGhVHoRX/6PnGEOX
JQQi1cCx1Z6dSP0cOLPFuyWhWMM9fLTDYK9RQQeqnoWbMj4QLOO4Bgrdr+RvqCcM
vhApK/4/Ba3vbE9ITGXSY0e8mApVzvX1q5InZM0wTaKUY7DDV8lyb8dEGGX9y9Dw
zbvCnjjL2I8Hh/RYX27xuuNrXm5ZzyU7ozcZALkX6VW7q7BLhECROR9kT6qCGBua
AgpGvPFT7AAM8v2SkWBCdESFmhLtOSupVfjeNTV6LecWmU1b4841pKMxXWMOkkdi
JRdbGgeUcwRBWUrp9kL11yxKfgvwgU//7aXE2rZCQ8/C1G2qoE2ijmOCO8AzIC3h
nXgrM1zQNtOWxcscziP5KRKfWdx0aeo8vQThiCEoPoWu8a6p1YR8e7sSqEL4D31g
GVh4mYyjeBI6AiYqpYkkPRAcEE14gxro4hp9L59m8pjxy/w3sQCN8FC6mVZI2yvW
ED+RxYq84fpTEXzceOcxSWZhUGMrA2TfV6cbsRMHxcJUw0SWjO/3PJj5SfzbS5Yo
28jKf61552bVMJQnxvM+xbmMTHEpRpVGq8gk0TBvQauxk8bLg1zMsjScJoYzgkGb
26/4JPEv/qTNEGwrP6OC/Rop1WpN2pENkNu5KWf9A1mQe0yIqtphUf7iohFTAv+4
7noMgAj/PxtUqtO8x7Yd6NHi/bjllfNQ8Y1vpvT+LtQdBWhExaJ72DkB6z74qx5+
znZ1u5Jv77S8W9gVJWiEQBRGSnYczf72fpnSZDhEKR4Xqlv3Pj8IWFLFuPSH6uIp
E1WwygtUph4eHS7uJuKdAwg4uw0M9G0FhdPn4eMpgRuhq4Fh5tXrW8nvlpboP+7m
2vR1pb4HHtqw1yRGMinz6WgAR2mC/Dw4Y8l2LQH+a8Cs8+iDzBj3e9fu4Kk1++MG
s6hR4GWOC03hFxThSipL1iR289Wcq2JkYwWOn+2Ijtigm+slAcw4zt0D9iG1tJ5s
iCQy8QexZZhMHw/1FK4Ma3YFRSRGQz1N/HA3HPW27ly9/uTujWevmxPZki0V4w1v
sl6ydL8sHRvjnet0MD/ZlCErDIGKMc7EEiTHNb2KGplg1Le0i6CxVkdNICbMCdf0
x6DnegolMP1G/aCl048rsnAFYIUMhg9OyyGZdzCmw+7QSslZd30NvMK5Zuf4E3ck
4d4TX/FG/4w9/kbxI1JxRkK7+s+fntUFq7rGRQEpYT1UFwiR3N6zoOBMbNC+qxKs
RZUsQlodHucaN6wPsqMN+vmvr0j4Zm6WAdOigZS4rjJdWzoi9YOy7H9yZ2OBYvl4
lyoXlgrea1qipUzN9uWivQTzw9cUIffbblN3ljUc+mFOdyibmOWsWShUJrr8+KDV
9nGnD/n3bLyniJcC0d6oZpSuHXpaFbRNPgtI/7XlMYAhnShY3YLsdKyH3cq+0tqV
My1NWVhCtiH3fzhanE9hxUbTx61jEbPht0Its71fzFRTJX+6/VeL8L0KZH+NTs65
qDDN92z0JDvHIsA8ans+NcF8I/CgHEouJEGSkno2J0R4Swh8N/LgDbPxKsbzu95c
4i9I3fzo7E1GJLm702IrI7kVhMqyj+WOtiKGQLNN8U0aljgnoMemOsLzHtK/TuBD
Lrny8cJR+nTmDEvI+07QmLWzFHDP74GfAEIRJ369yNLPvC+HQfKO/fsxvvG3jCqD
mRVeZPkCdbsrWCjt7WwotHcMZ+BtbO4L2Gdyi3113U/6dNSnc1mvjqOa2RoXeyY2
3zWbLxqfy92WWPHwfPag7vYgdQA8e6w1pa6ng1k3GoAxNyY4SW2WCoBa+pg0dm5a
jVwf7s9shoKhWpfC6Tw8m22/7rCuD5tECd0wKkQz+tELbKbeYtANc6mUPG2azSS+
K5iitgnTZvM4PrgzJon751J/+4r7KL4ND44qHoWa5JyIRqyqngxkeK5ristDfYKf
OLglAK9C5L1cnn0BJYtd5C25bjSdex2U/+tzkjD5jGRQ0N5MoQLHQX4dKqFX46at
VTs/H8xbgnvQrpDm7uvTYkXJu4/xMxpGqtIiPuMPjXXnaX3seSiRII/wZh5O3wk8
nJQuCjK/+4WZd2VHYl3JDHHyUYwX8Ht6oFLfe707EF8oCcLUfd6n/Drh/+FvoF9n
X0o4mTXDwhgL0uIR8wFBCzpDTbBttC/gsjUPXu1zlxln4XBOfEjaJg6OVh608T8f
OLYwNNLhZdakFgi9uUPfS8VBrExX4LtDJtYcj0yRDeOnySk8FPWHHsFUbFLlE8f/
8Ff6PvyxUXxfXqaMT7xnaw19cVp722tp9ALRnT2c+l1M8Y2a5N+mIOVlRvCUuVmk
R94qJvKXhkfQ+ijHn4DS6OuOgkvSnfKwBHjThGKMM8hofpU6Tp6YyAPnbqdiMfVy
j+ippqFbGkaUdo8EDYhYty3a8AeCj+2ETwYVoZLfnF1d5vnTxrDYD6FoQC+MRAJH
Ka4FJHIuUpHkhmr8ZBjrwmENNSt+vUFyb8kTo+JsUOOPVD+mx46lalre4HebOZzL
wJ2D3U92ELkwjyTrElcRzP0+PgWY/ofXWBXgx0BzgaXZzYSBmVagOgZBIslZrzQE
BM11GojNOoSWNbenBkwG8s3xMETi/BsePE7e243zB7VeLsBUn2fEQYG9V5zZw4uW
wIxDDQWcWymDoEaaTRzI3B6F8gX9hxhIKC2QgP+YjjupOi2dlxtSpW5sqBHwadLQ
JlxonqENb0KLsk0B4DG8dQN6OFt0SLGsbjSbk7EVEU4lmYjIkLGX+uTRO0mRXRXs
lAiagUJEdzX8BeHCqgQboNt9rTGB15WGIuKQLPZAMAfaLQMUhKo1vozwWhL1HrfX
WLibL7ckAQ6a68GkzReEE/Hux4BKlv8a75Do9U7olly85eE5C3ewBc7UecYvxMaP
RGSKzHbhpzFHbrKk2xyjex6XX8tDzxDUco/JEoI8+Qqc/Kd2oYRW/m/d/epw8/OM
dyU8ZmSgv9AisDn6SOEBF/xZrAeqGsEVfPSVL/7JV6/IJLe4qauRz3y7ij5c1Lce
qvWltkK4pAZXPN8/0tDCZxt2WPCryBMp419oBW78sYKMVC7axHJV1JM1NwPdp+sh
UeE+qO4E4kpKAWBbBIrk3D3dnPFmXEyfEU+Tye3oXMxMdotQ7w3Z7SVnzSfn7xiK
GjQOy59LJNLkzUf4rvisBAPXF/BSzaK8H2pLK5IIEqPK83leLJ35hOdx3fYNB0n8
Ynii49CMNZLwi9l52Hqex7nKzlJfB04rJ75otjg5fCtCN/d+B6iHHbsUpi+OljAJ
nQLlRdKM4tjpV3XZGN/syy62fFuv4MYKpRdmHn3dsNbi6EcT7yzZjL5V4C5YIjed
Rc36zwzvdhLB2gXl9e/0s5eatNMVvfIBb7M/iV5ld2wpKwm9geQbCNN8LHumjG8S
+XjgrsB0Anprs8MAEwnViC5rV9TrcZYfyBIGqOi7+kBeSRq5opC3n5FeYqmfkeX4
6r8RBUsQtPN55o5xWNQpKTmsBVUfxsN/1Kq4+VbEfYxjibBZimg1sMFmWBAGw1ie
6MQW8BayxiSLkrYk5Sb78itr7sm3rN4uulpsOJeqz9aBi4UzmPbdI5fktcyywiYf
pJKzQKENjUBPqqoH8RG3ccLP4+IzNDAkybgOAWva2PmINBdnTPYz9Ih5t5+0YLFz
oLQZHbrvlgPD1MW+TExXoBVrvARaF1gjlOT1HCTt9n3jMsSjEDrsSBKz9dEEYXAa
kV9f9mYIi2D3evn+TJh2fxVfghKZZGdUEZTCWeueJQJrgSBBvGEGi1lOqRj/DrCV
M/k7e4t0eLHOsZtWmfmPnm0ssek1pAVrsJuPy6RM9+2CrRgqW84uab8yxQfC0pBe
47yu1aYBEB8K3lvCU1WXHDXu7wgd4msZ03iso6k75oMm8HbdRtdFpn1EnP/Y12//
xLK4QU6XNWSI2EZ9QjhA0f0pRSc4yjOa5E3F2AvPsaPr7EYUZJL8RkIDeOgSzp5X
ah03PYORV2dpmiHAZ+Ta8A5aLTDq/4j0DCflurPGRQ4naUFD6IHs/GJppZrUqeZJ
LumIMj6mMLSCu3To0WyUs2PwZpMwUqbzpggw2flHNQkYFSDUpX1z3ifxl/zuj/8l
PHqAv9G2UTLMRTtbj48wfXgMnO4pmhF4BSj0Se9SdJkwJXqvxaTcKE4uo+6kL8o7
JoZyDVBBibO4OFIDm8zn7x/bH1DqK/vT2fQbaeLjC/cUtPZXnPolzb+ncAQVYfL+
2rdsWFOrnecLp5Yge72micj8ixmuOW5aoRyedxPMqHrrtia9GpUHB2U2louUtvFb
ywy8DcqKWJeb2u0e3jSZw0DaUiNsOMkcAzR2+dJVUXwnd9EMZtBx+aBlfG3AJVci
+UKM1K8nCLKEuihCfKS3F25vBag/cXeQ5TRgv9anRfqPK9FUAv0UgzdNrzTmJE0T
gJhhQGrN6SD/D4vkXqiX2eondpUuqQJIPKfh7t1+4xgRj+2Cgyz1/2Yat5NB39TG
DXhNZ/OlzJXdPpffxRJRu3Q5lbOXX2/aGik7J8S0+VkjV1LEN4dqadOI0E7FYasr
q1vwvfjrDkAVPyvrUuMifndsqx6PPvJpWRmDFJ2lLRfapt+LZ/+Uyl9l5XkvcZ99
CcUprQrk99yzcZgRj8lGEaGlxyxjPKZPR5LMi8Aj+4i+DJxEwL22fC7X8Y4sncex
9DaGS3HZjw0CHzGTrvbGx0O8xcsd97/Z8ClNjAGVLn8Q1WHVinSL0pg1U9Vo3GDu
KlcIvLe7m2crAQ6eAyZAhnUY1sfgKeeETh4wsoQ83WD1ZlHQxS5RY+sbONktHnQa
aWQUOiEK8EMdW4wLQzgm+WHvaqTttysnxyM3QZfhKYtftObwCK22IZqKfHpqg1XX
fInfESLbVh4GIda2klPVq5gIiX1nVZw/0Ff+v5sizm9L10HJDMUkb3qb4pDRjiRq
k48EhwgRUtUZbkAvTVTjk7DBw5hZf37eU9I1/nxsAgqFvfZkn9U/zb6UQr81xady
COU6y4bw1A1teQnNSrkqXZjlrH9AXp6q8MErxgeohMAbZKNOKXl+/Rr5RPOppuyX
ih/xZpAh3zPG4JHGlMB8lUDdrZdvryDf4DwA3x0NQP7CkAbuSep/J1zalQ8+4otu
LusTR1U8kIvw9esT8RsMeJU27MDgY+FujZKQE6HW6vgojXjRVoQrhGIqAldC9dQf
U3eZaNqa6ypgYmwTm1I5nduutnDHnGI4lhpo77g2lCQocQuLOh9T0MA1RgtfwRhE
mRrAUdfBbG6nJGjLD4DEi0wIvHcT3RyOQU2Zq/W4UHfdW8PsEGAJ8oZzJFEgsfRm
a9KOnxQpzcfQCv40OXU5YJbs9sHuAwF9zDDZjdD9Pl8U3K52XelOBUv/elN97sY8
+guR7t5uM2f54cK2WI9WRGVyX9W2FOL5UxGpcNfAJwDUkzkArSDux8GzKwmuXZwp
tvmqzLqBoem/mz7XaUOZZaBJN6e4Q81O/ELqsVUt9wHykwsVMwkEbqDeFxXgkvD2
wHM5+GjcDryadQYQa2wJErqubQBbuoFWLSpSeQBksvwstH/h52Ly7+DCAm0j+C9g
5o2i7b/bPX/pKW14rDg4wIfIuwI1p01yyGYU5PoNjPOyUhn+Un6pplC379M5YBE1
XNR1JH6BMsiSjshv9gT1YAndKpiF6Vs5o7SaoQd8vpT+SMTengL7uvHo3HIe0XLa
Ou31vrtk2L7yXH9u+YBDri5dsIvgraDLjN3G9ynwPQgAQFEEEDfFSGAdBwD24ISa
OA+op3IlCaGXmWnAevgY+j7KiQdC377poIwbZHCpjdG8h0u9ABGnGL+j6i9+lWGC
S4hU8V3PM6dRcm4wT0rlC8w5ioFOpIvOQSzktsAtBrdT3g7uZy2fbCu1l5KYY1B4
hkM7hkFXYgGDJxbtazox86DSh33Bh8ENaCPrw2AEu+tMfVmtmLXf2irXAQ6iXMOo
n+UdbMEHOB8MV4+G02mjYGbybTOYgCE6Zw7ETR6J1+hpov5gZ76rGGqgUt3oKeDg
kZEwT9a5UsA2DYBVYp0TTTJyo3+6ZDTdF/Z8i1IINfi6bDeWD1TW6tduh7YAUTjK
nvKj9Paj2kbMESvkAacE/J16HrUkbV8LSfVOnkFeDs4Vaun4Cw4rxAkq5acAgwnk
VybQvjfKMuG3TYcbRhwixz2XpvV9fAWsN9GWXrFlJSgESY++0G9Zn8K6voEHXIEK
FtLMUmB4uAS7K9TmNY/j4b18gKOrdjI3CZfIX70AXD0w3+ksN/KJ+7sx3VYLsuxO
NLPIiKcn6VCywQoHQg7VaoTUqiAp+Xz9rlxeEyZMT+9H8R7stua1gr1j7LdEGfKU
Ow9sQ3WABEyXLZgzEgHZZOrlae8t9bf8wLoLod2LQqlHMisr7fusKGLuuGlChS7N
JrqMelE0f3FjyuKV9Dkfgk/QTQP2aZHUqHcbypLjSPxEP0LJafq1qQwtFhVioFg9
fVANGQt/UMbHkfJGgQoW9nmKTXk3PDx5vv8PaF+UpUprC+tT7FoA7N4pKh6oiK/X
rzFQi05ZILUOb9cSzG4VKoas6w0UBIl+q9xQ57Zj+AMaDiLWv2r+YftuhTs7dSb3
IkH/S9J55rHf0dpwpOK+tx3sRB2mERRpsktcd+ky+ErP+cak/wGec4kU5KT80oNV
8IOXt5PfCMVFpnC9f1PFGeEhWD41klogCWijqqRQMHyBemIWKvSLHk1WjBSqsgRk
llMKjjc9cKcfW98PoxEH9jf6PXTUyq7ixep4++6kEOncnTW3S9IEYDZNZL8tS6Uk
Je6dnV0swcjC4Vwx88OGB4Z1KsTTeGdGDuQD4Dz8NTU9ERGtyQPj20MGRcaTuT5r
hmmhUjtP0J27UvcnqXyLp6tXU4jqBLzVCBPfZjTNvonve8Img3zZDylPMSnq2+sD
yICYilCVN0YZOgSGNkFB4dlP4hCFM0dfCYKEmhZjp15Hwk8r/LMv7sAQq83onW5u
1XrKTo5ZGGnnO/iisdtkJOL3NKYMNytfDcsy4HPvZGmhjO/xDUwVaQ6R0noW/q43
czwT/eOIJxpnRHZWqP14PlLvi5hPfq2T85X75GG4aOxk00XaEmIlHIJqPF9kgfK2
/FB/Bqdl6V+3KcY3Km67f6QlenTrhKEFmM/tpAk5nEPZTDcm8/KSD09aXR9aVSuq
iWo7MluMHjLUTxdcABxYFy/XAOgCRUMVhwnSuPKLe+9bgdoWqKIauXFGeeHm+w67
BH+OcPanxSjhC+qN1KPu2YgasHcMfXEsA5Ywd6ckxoPrfZzoX+h3YlSYEyP8jUr6
lizX946/jzqayJGPVmbX+wL77IVWaDFWkuFTCndxml0512uUJwUcsmF4rq07MncP
fvan89fKfAXX9aZBHmBAKsUncJFskb+AmfqVMli6Rc46SBkvHR/+z/HRXjt6f74/
hXSp7OygPgW9Ub1Kg3TMi+w8wZm6Dcsx/aeInE+Ls6FznPust/dtBkRXZW/vizd9
orjpMdLTQzlQ3YUtQ/vgOH4SI4VNmPBgVgaQNDgn3XXzRiR9/zCVG8cEO1le74ZT
pFk7VgibaJbUsgYz0wuPxkKKhWjr7Q1k15Ag4fqUvxJTnOdXC7D4em8opybjUpNN
ZWvJDhC6oVnnA/9CHpuAwlg6jTjmRY1PefTIcxrRMHaAsjSEuvD9gcAwQ9MmfY2z
z0WDQv+IRK/vSrqHEqpV7zTfysQreJGY45X+vDNhZWvD9a4mR//IR2HJLs61J3qS
l3ylYXNyTm/PyV7xaPIYPbfz2GgopAez4mFiivs7TXR5iNPIrWp+BXSkydp5/1VV
U3hunL/J/ohVG6hw0rJs149xC8qaHj1haI6RPJaVuLUBIUO1O4MVKgsd94DBTBdA
Nm868F8HcbsROcTNBfEZhsiytQQmltqFq/7S07UMwO3w7u2Dqoij0nTlUbMJqS94
VRBgmymrduw/4VnAhM1TBZDqwRGl7XaNUZBGiDYCy7LM/P9pD+Y02wFGim78d60e
/pUT2ID8sgZDtsYPZrFC2k8rssjq6KpZNDqqxdsbWrW6wfH/ir8cpPOAeNUvQl+b
IIpOHz2rQxGG+JeG1aJJ3yai1YIv9L9ZvZy5hnvD4zi9mfSmio8fW/RiC04HRq/6
92MFtaHeLuDf+KjmwegVxeSaPY5TcBwlUxlXbTXmMehWahSQjKy/JrpT1a+O4hJa
DZNuOQqOe4yABn0Vtaa7a9bplfFxi6SUziBz+am9+LVTepCrMSPjw1mmIdknxD6U
uI4ZNVUCUSFJEPHUKzzlM0n7uriMalmctoYEdLjHztetfqWJia2W7bH2/JHqSb7g
t6a6k7F1j9IT3y3xp3jLbU7rJ+YqmPsJmhJzZqz3H4YgwhBE9a+/quS+enPJ2PfV
cwz/PkdFBOADvUPoe5buIqKsmhuKS5hpfc9jndKn9XipMgmyM2Mf+WHotmiRzFyy
nkLcYPjgetYxIbQZBTZYXdqvmm3QEQ/mw9p/IjywMcXSJKkeYCy3wz47An3zPWut
h8gJQ7HRCbMxSa3TB+hxqxjqXI1HzIY8g+D54+tCA1yukMPyMELrZIHQlWy+eVLx
EDwsjI8TQVMjZwZ4g+75mzSb9buimFUjoY6x5LDkwCZtpCOxeZwzTJXkCiqU6lg1
dnHH2mLWpZl68zeNw4jQWHpQ1xblQjocaJsm/DpyAGx4VJ67Iptmj0GEvQYGgSsn
+o7y4Cz4FAzUGwcwO/ciEXhpOo6iFL32ppIN8JLjbZrjFw27biTWwMENjv81NbjY
AWC7ACcyrRKBA+mMfhoV0HTD7WqXmlKZuZHgGTTafsfxVdiYQMft8LcWqT/RPUTw
zVPf+Exuz4BMmTUsLskSR814DfsHE3kfRJrMUi0CmcpfDCuow0RI66tIMSE6nixb
+bCeuy8FHgSgnIFJF0KPBtrpVNppqfRa0UX8Xak+gJg1aJZFnOfiMVA1DtWypRNN
v5QLGhK/dir1Rf900oL4ewZLdZap0wOyEFWuQB0GyewnPcADWIzYbGCmcy16CqDU
poDM7nyri6XbdyzMo0kXyJ9AFXVvTScjL+9BAHGPFPTyhIIXohlJDysNWOIo/3S7
hqdM+Bmng+m5p4EEoKFjx1d3Y4TxNRWoF5onqzRwSEj+z7EdkhvD5JMtauLVvJBd
80Pcuy4t9s+e8f6rKacAXFZUHgJzUN50FV8cgKeQx/drB5XtEJ20+jmGJ3kT60O5
Xkjax0qi/3kboWv0G6bj4eSRRnb6RLQKLTAu1vcHVjKOUgpDfQqNXFVLdeJkMr3k
mnvh+6OfJmmb57NZgici2OWorB0uvwT9sxU/bv4mrKPgQaQF+gz/Ua1W2wAB07CQ
SQnffjic4NxoYOD91HMZdxzc6h7h59Gb1Od0d6cFEyUBWCB+OuwEt1KwlIjTO6ko
KtPWYTQU8JH44ZLSpwfv4cXAnJdt2/B1d1BwaCYuHgxfAksIbQA/ZWgMTIDLHEmi
jxEwcwned14DjOAosNbsp7rZELiy1g1IJ6aHlcpz7pZDjKV2g4lq8xK4by8Cv3hd
dCcYBPLbXlo75DoCYEfdHM6nWZZay/4oFoQSdxVmsvMqDDgXj3hF6h6A3L5cpsBj
a/CovL53ryoRzzaztZwmX7+ELcfWQo4KgeAsil9ekMyk80TeQJGv2A7yfv2Wo4ZM
EvS7/GMWOmeLnCstvwvrmbqQvVAUOsD2SBQJsFQPP3Wp4ooV2vyo5+qOhSGpP8th
eXw/D2cgf9wdRbMETuOp8fPZ5+mbN9jWZGpGoorHwp95oTPqTtD78RnLhLSrpjU1
cc+A9+SXmxa9GcRDJ1X0rGZj8msHaalMjeGcSGPugYpD9qHmtbC8654iFNZo0fLI
LtrlRm7vQ6juZkNm8fLVGx8lJFLRIHl4xY1n+zXQA3sb+Q+RamBxz3/J0OMbvCeo
tBZSGbMDoRACpEF4H3LQ+K/COT7Cl6d379JsSwYRjjM8RoZos7+gi1bPMTG/1bH7
QA7u8rwVKfJ7qF9ncjTAFTBvr76Hs2GPKW6Tjx9D5V5SIudqv2cg8Az3S1xaDY2/
S6jy2DIunUw8JiU0PAKWi5bRI/J8qqYEP/e+exnzAs+loS3458QhqPb3Z/cXM708
Q1YXdgS4U9IdgEIyQ6Vh0U2RU6waN0b80SzOPLqdAAb9gm9mPqXT67V7Le1aojBL
+1VLLd/2P0HMnYmFU7OvktvD0cywBW1IWvWv7ZjorKb7VsokKIwhFftpXvtSS8Do
c9HQPKWmk0kUyjDLeO0YLA4X4188zZ7aC2rml6+XTFrMyQ1YKUB9IpVYqgdyD8Iv
oDHqVETP6w6HdrC/aITAcyNq1guyTQcXFgnDLaM2/0ZCMEXKKeqz294LdT+m/lMB
e54GMGw7JR6oWmoFKTWWZCoLR1582gnJr3PUzV3Von1hP4pTzFXN07kdwv3gQtOG
O1zidjwuglkPYoSX+Bqte8EuA/y/0F84RIwYH8EUoT9q5T7hsFYfZacj7VWwf5Wd
VZYxitPrnsSRVFEKLEv+2+o1XZaqdaK5BCw/ASiw+qtGkNwx/yZIlPiEP5K1YySF
nwtFDfZlQ7aJIE4GdkkpFrD7Aki3WiYs6W3qAEEFe4tdjpoN8a4FMDvdflDx+QHv
6HdnT44W2f1U9Kp8xrn28GpwoxkGb5Dl+iPZxdssAz031nBO2M8FWhv0s9f1OpUh
MtmqulYDCFKDmFbvOvl1++BWt5YGe9nbszGd6zwQ5qH7iCrwDQ68SqVK2qJk2yIZ
t9gpFdN18l6dAFODb9NuuZeJt8np1pxnBCOM/FfUJxxwCOnjYp0kpP2gL1KoCbRz
GuwpTZ/2SN7QmMR5ZJ3TBlwp9VjMERl3uJn0x/tMiPwrcK2UnlbATxlLfBCBDpME
tTA0el1X02A8XC3SoMZvMLwuCK01pZ4maCrV3z0wOsBORTH9ojH8Vkz22933/BMW
ttp7bjJlgRlPwXoki0M9nXFQDu+46mcgfpSb009evse7Z5Gb3rtGZj1ok/rGjMHn
CB9qeS9ouj9WnDEplB8gWlZtbN113FqG6w4WdHreGhFi0AQRo5Dx9ZwyQ3I4tB0O
rsmWXA4MJaF6VJRoZw7jLqkABR3anek/nc4/ZmLNYot7AcQGCZLE1cYZ7MRHdLA8
MG5LZuDUcY2G2tlcqI8COSLYlDims5pPb6vnhqoaUi3sGXVnlGnEWhTiPObLDPEO
5H605Md31SNrTjC4tcl32SnvkBu7XYnxqnLm0JrHZmYLgzOiqbFRgy6nbqNmtGSy
rKVDfQsB361I9yKflHdxU1lHVxEej2wmeLf8UcR24owyRD3Wu4TpivFAG0n5qb+1
0BlLyB/s1rm7FmjDbLbmTpJGz8s/Db+XyI60pWRwJFhwaF/IL3vlpQDGm74XiyWx
uWLvSRtRqjDk4XGuYkUyQNKboFzqc8KZvcYm42Vj0TXFgxDQVPKk628IFbNMhJyN
ulK/oDg4qaWZOihF23kDHqK48qB8ScMSc3jYdSq+c6ewEnTijGzcUNikS+WlXpT9
Kew9vjC7oIVnlvRt3hA9W+YQgLgRVq8dFTZRZNOc0sQCqkIiAT4ISvOWyN+06EVw
gBpW2Hk1/s+jpydmhkPKrQEGgWxJhBzy5wDdzIOgcvS+DFDyz2X2YlRnzLev6ckO
UMg9841bZruVcjDxAh1NbQ2Y2AOOoxFgZvDVDrlxVbDBjPAb15uamQ8aX/l9i41S
xJJ/w2lmezBYHxtGi30pIz59lMREvkQumdJwOzIr0BT6kMYEIS2x6kszzCkejPzk
qsIBR+2dc76kduOzmcpAK2iYWj9FNewrGnTfptAremau0w7VUcjcbQMhWir12Xau
XPtOdzJ03E/ZUaGxNfrl6Qm3cisMwye4dRJkqyuq/GRdLrcn8JddwMAbg/tVcrCC
OTDe5zAUbk4TSprXUt3mUoq3h9TqOm4Mq5Pb+tUYbVCwakE/12rAkAooNhN+1siF
g9RLC3G9+cDys2Ai/x0yqxPDmr42RCQUvTD86QW559cC1VPXOhyq/YtnTfCZ1QCs
l4evThV25om5ZH9rYa9rSmZZ7tFydeQI1NaN0evFKTj4KFaagS3r/K6nxawmn9Yv
4Z1E9uccXrI0tQ4gurvOAoTUsyy+9hDaAb0IKNKt4nBRT1R3wpqEtYg84yKQwTrQ
8LFiWaoJFSyIpiliiSCoxqyt5LfL1xio72DO+ckiWNN3u1WBkU0quMhRXj7DYFCB
kP2/SKUXajsUxblkF3yTwpgLOKy5gS9fAyUJZRgkEjjq8z+sBrS/yDhjZ5hzOl9S
o2V/ZFc3nBirIk1HMWlfxVnkbfTj+jAqa2SCr1GL6IXrWrIuNvbo0soZ37gO8MyE
WrzAiLlnBkgbT3qq6yHNPiaMgGnC99LuK6GXkOYu8Dd+Erk40CklI614IC49XHSC
l76dUFjU5QfFAgrhKDlRfmY0G4d5mSabIUBZ/ksL87nHQdJ6Ot/lSFj4yZt9I+v1
c1IpuC6yXVLeZyZv/qfywPC5n6lS1+qNbEMjJZ90M7LOayLYZ5dqC9lLMf3XVbWd
peOKjoCMaeemfbzZExUJhcUTQJ0tFH7EgZAVUm1K6Eu2KLlvRXqDBrlVe/VpsEJu
RdsrpawGgltYL4u6d3TwyZ/EyNPFvrf15CXq4GpT8LHJ3BcUMCxsuErI/I2x/Hqf
b576lolFromEG3Rt8CcBoWKkaEGycZ3VtZGBOrm+QGj6jVWhftAFYhJLJXzjHV3Q
N67nFV9myRDOSE9vA6j5OPwInz4FQiwzSIoYKbLx+mWcNp4M56fwJG9YuJj8XhNi
chtP5He21rLTQwozvfYy3/v9iAZ7XWwUdBD83bniIhl6ZKRKVXEO9Jwu+iM5vkCy
tsg+gapSY3a2KkWf7zQfjLufJT2mIRSFm3oi5rP7ivB5tzJvvm5T71cFLMjC7cic
uz/wQqFAsrkRmvcNZft5aDe+pa14K9D6a4x75nXiZIcTk+1qehHLzQp17AfhVkZw
tPsPjjhJnLMsHneC4Ld104I0tRpih1YcS5iu/V3t2/EO9ddABlABFgwTx+WvM5sq
kc+lB1vDM0SVtnd6GdpJD6Etk1y44p1s5oab3ZcNg7M87Fx6kLY9orKnubitRbJg
PmKBAmH2IoyXLu+nyMJBalDcf7ooDNcRJYBe0b19Efo4rtieOZPIPtnU2Vy1hGNX
kJALQ0rkJ4pX8GD5ny0tbQ27ygwWYDZjB//LJ3xdbDIOHVQRhOJE+1LJVbpoWh8E
ckl+R64Qr/8pTTRa4Xpwpm/Yw9EFlglSHWv0ri+mdO3JarBUam5loYWdO7vf1YTG
Yki1okYib/4dO0/zu1CIJtOVPwLzuYzz9WebHzkO/oQPvi30S1Qjf7LN6A6bfkqR
mdyjd919WYgozWTjfKhZxXBp+27CUKTAKrvSz5fQCdq7tdFNRgFrK9UzLIWFdsnA
b1gSQthcLA+VofEXf9EYkb9Rt0dGQBvJghf+/ZnPj755r2HL5ebsvpV9/GS3BOgc
vxxt7ge4ZAqweaVVOCbIgTsYUfc1DQscqTInculmFhR7aC9pYu7/dTWqItSMPY8s
9Z9Iew+kpU9nlhbCF+3MbjRVoVvv5CrWSVP6KMdczCWdvKjQ8e3UKZaM64RFhGA/
mvUNdYz2WtuBwEzNt3WLy64NaNuUa+LL59uVdjEWFusnrT2kik9Yqsjui8hfZD4X
SI9w1AFYDsFvDzQn0CZPOSHdRhnn2yoUPhHPTQW5w5epcxUGMPiIDiTTqXg6eCgA
PU1oqkjWfUsJfHNJfXwmy2u6la8yPOiX9eK/t02FA8+phQiPdxiCdq8rZhrpR0BA
XncSrb5b8nLA4/fZ9NO0jXp9e2xeEmXDyFfIqElXrniFigaJyzgpQYjbrtVjs+wI
wsgOwOKtEJ+fEE5lxkZzxh8P5D7RQxAMJLUPiYTZIGRgUJ8lZSVmMhipufWOz1ik
cbN4Jx9KrPY0AUcWFBXi8WfymIRGhZPvO2ZfCyzQf7uKETmRlEtHV+cK/i15wlJS
5BatbicrgYwCAjsxfBkADjutFdYtLiWEbTVfh81r/S2OE38mzdvSJ7aZnWzKNmoF
00IYVDct5eXokgSTx3opgkHM8dBASouTXRi5KDm4mDrK2PqgQz8xVJZmm/lqhlix
/InKasHSjhvWYOR0TPVCuPxxRkbUSweYMPs9xd0f3vB+QsMiVv6K6UHD9/6I5KQe
eU3JIr/akPa1tzb7ojoxVqfuoQAdMXFJeb4NOfNYF0KKzkPJMTxBkmE8DVgkEhVX
vU6fv74DpodKVtYE3F0bc6SV6UQLX170WADcOioIb80UfQhGld1sMC26oy/363mm
zRhKu51sGU24M4NI4GtDSuXE35b0cnrLP3BkVNE9/2BLsAZ741MwGaCmNHzDeT1l
RZ1EtehHGLKMXgoB71UU+oq1gQx3Dk84PcMgWnw2ChvcTFQbfbaDfojlNZ3GxbAl
93I5MB/P9R6Dfl3ie6qXSLyjo0I+eX8t93EIbDi0slALNYsRhxNepE62M36RjwIF
UAAV89BHZHDffBYrGKLAuI3hGDe29fEdLHAN7DnnD3kqiYWaq+kdEscdIGkDUBul
ux83Nmf8So4xtUAsVcECFglHzXkTpp6aPBGWI/8MRo7XVtatVSSV1eT93ExAzsOr
LyXee4Lw4yZCw3XOy6jOxoVtYiDUmLfGlXDTnHyh3MJsgWBUrWn/+M9cE4TZn58A
6wocka1sSrBAPHnmi2XDcgT3A0YFApFJkFpWr2ZS5+R3+7/6LKxd6fXY2UtuOpaR
nKtEVbFz5T9tWNznPsWnJpcugxBOU+spS7WSDol/38GU/8Mm8Qt8p20Up/RVTXTH
E+a/WxpV3ioO6YOIUzUuI192vCY4UbiDGlyoc6I+jrXvm6mKNmhF7dVJpUZEipkV
cFv0uIk0stU3V278sB1PkqI98lEBQI7EiAsBEBXEGG9xCsv1scfu+eJmdtl1ijqO
ylcJwXczfQQsKIDsJ+73JgA/oEqUYtUoWOMpjT+dzUlFqB7CC8EUnspK2QlvOGNS
VHC6vLfNsbjouJu0crcRmlHviSPZlaI3rQmNRl4t9OtqykiIsQ2lXUDr86/Noo3J
ijq3k09UzwzwXrjXga5hIMAmeNu+hHyPyWP8bfbgFKn5zTdCeEddD8Hk19vcdQPE
+6zcXKdaiagrnaNfTPCUqrd/Fk2cBPHUC65TobDW4V1ulypEkVRzDvnsvsxj86Gr
1hrrKJQ3DMKJArRkE8XHmTjnET07v0usWvGBrjuuKS5zx9HakLDWYXPXK/T5UoIi
H3VC2u+D0g0i4gSsdONbrvfwNcJVy1uPbax0KHRfSTqvd4tB77DtYIFsfoaS3XAt
3cHlPDpXPtCaZAy8bxZLo2zUvL6nbiDxHmHYfU4kAbK0Sz3J8Y0vuoS9CNq5leLP
KJSNpKhxV4YQzHmJoEuLVPG4F92AlSZBa/wYBPiwgHsL9riMzTkwJwZd7hvvYwTs
qp6+XZS1ZNnfMsNvu/fnRMEuje4+/VHEsvu2FbnrFoym34vUJWjg+CfHYGbDRi5E
9y18xfnb8Fba296uWYpiC1QzACrZgdQyEIur/cSKdU7PInam9+CeoVT3/3FtEepx
7imOdCF6z1LxyuzoneleLsQaSIJK8tdbRzNesQ2ViJjoY0pLr2K7bCClL2eySmwI
9Qv8sDYHQlsCiYRPl0zO6aQEElk3FJY1Pdpq2uO46slBokFKlBEOZjGV59bRi07k
L+kcqk/8ZO2nrdreAQGGXSPmqvwEw+3UsyjhgX1gc4KG6cLN9t2rlC6qngllyHB8
Hs4mZ0aWW+sWFdQF7r+cP9tSST5TvnSAXzrm5lVRFM1U6S/qbspt8bFIXFwHo32G
fZd9St5PYEgVbOVf4kFnQc3cUVNRPtLvcSmYVTdX/hXjQKjQvw5A13clGabSm0xj
cmE0P6ib+1Knnguhki9Vo9rnTzmVr0q0mPx1XkeJl3AJK3g3y1WcM/u5iBI+ncbM
UqAPyojZarB7IH+PklwbPciC1SdyX0Ajj5LZlTtDM2/StBZxnnF8dEf2bHRhEzFP
peVycgoEbhiChzIW8cGoZJAJdEXVgG1zpYwfjfxogrHeo7QFgRIxJKp7c5LabTAy
UzeMArNb4QiEwL5mcdLchYx6ttr/drSAYgRvpWT9/K8I7xRJGf4EbbZoLlyvUeA6
LQGLm/78KKLT9b8EuzLtVkyYS+MfkGp53QlzIuY2TtXFMwQZviod7nZStaw+/9XU
zIzV00HRtR5QRn3LOkk7pIa3vS3+4QNWgcGqfkASaQftHhkMal9m6E5aHIEmvUgn
exR8TGwyM4qO+H+VEhjwPZZa8nSe5pj67PkXb1FwSrmkeK1jRfT7XSbWxg2X0jv0
xebCrhS7Kpd2WUes4jIqT64e9LOFNTcm/K0rbC97ieDxZVQGGq93rudzGGljepYO
uR03zQEGnC/sLYnFB/N9v3M8G2/ALHZ5NOtIo+923vlzHIfuJOdMpD3wsRca6oId
xA3NCCbgizcSzyRJ28HyOGKBWnJC1CcJeYKwliHUoiy9AqOV0RkGJ5ZPtpnZ0XrY
mxzLKe2vlQrhCvzNGlX/dKVjpKj3LNQfe7rO2RHdR8JEoc9reqfvV7gAoPFlVpA4
3IqkdOtrIdijRUXyrS9ci4eILhKFCVGEA24sj81QkqThqaNBYEVuf6cvXiEnzQRL
q/piyfp5Z9qsJdrfF7HE/NGAPAEc3F6DCJhxNBivW2cnNa2m0cVRgX4wPnfYJMiX
mgNTNdPImz/bRLYcmx+swoC6lS9XwOruIcvMlfIJpa74MfrppbLRY2y9WVHAlPW4
HU/s3WcDz7Wz30VfsNpFqLrCvblf9/E9v8WJo0+qiYzQheyjJSrhqDmzJWBRucAv
UXVpzEJbfc1vdN9w5vmJGV1FPk5xGBiNl2gHRuCqUIL9qsKV/XvJYaqckuOz0MWm
`pragma protect end_protected
