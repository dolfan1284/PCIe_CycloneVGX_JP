// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:56 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f+zmOiZ2vprZ4mfRLFVagE2t3wqEN9slvh3rgLS9qNKCxL0Oi0Aa+HWYievcIiHh
e2/mtwHptypyYjEtdbXKr3lPy/IoE89lIhGjMSp1VYzP3Nu/hF22OGT/5QyvzC5T
fWQY8Be11AE8GWWreDYqJIefMOGv63DGs3jdJ5JzGcY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26032)
V8YIpxG8fDSwGgKSUW6H3PiNXNN7GUg8KOFk7ieKFgdeottyICA6R64l/1XBpGHU
1PCAynB04XeixKHkN6GdIAwAUH2okBHt+MAdWGAsW1dR12oS+4fIICb65GTCumFz
bt/FbcTxK8NLBwhEUgImeGc1zg9L9IIJSwgj0H/24UlVkyPnqH9MemtJuetzdegv
DI/ZCumAm2OJaCXh6VRQ7pz9RJFCMEi4loG3RmmGHaoNbr3xHCUnrVNiToWgE2OB
eIWMzs3H4KoAhvHVuE603AtjSZEfmNVbu/uq3JV1ms7NEpeqwXt6z1KEoikzpc5Q
egyv3+x8QSi6XcMTtYcxU3I8RnU6A2lsC8qWc9AIEHvHE1QVO/LaAh1L2NEmWjV5
7WXwBkyiO8IZphxORYFO7j2ypixI8024M2LsqghsU7BjUca6WsinIOrTB5fCyjpu
H2Macsfm1w5+zPPumIGsB8DtWn+ycR6G4ldB/ja0sp6ZF/qP0vYi9a195N18WVKE
DGHc7hSyZyYdkOSBtgnICINiNjaxHp7mrIjLABzPzMmWNxoW2lsdoRppvtggM1VT
q9O5/9Uu7H4uR08TnncNc8KYzgGq4CJY+3fzjPYWj0VbXdU02oJ1KGSgpmpw/Gga
c1vi2zjlYJptTINbd22NhaxPLu31o4GhX1bUyRlRwSJ+yqTy9URd38tNubrVPVLj
KE8ELqMbBFQ3maSFnhXRAhV908DIgwrX6kzCmxgAnhAcjuTJD39YVmdYZtBwByJg
ccgl3Zz65+x4mzIM6z9O5IdLmjX1CnK43aDL3VG/d8/Dfb/KchqNPx1h4C6Nuv2w
BZyTZPdHM4xKz4ZvGTRV1dkfcYSBWGKksRcDYR3r80wE9mhrQnSs0LEHLC1jRu73
sXC2z/5wezuQo7kAAvFeVK1cU15dBYfQOOURbpu9poK65IcTts7V9RQGY/ePLKRQ
wuuZlqfy3VVOcVcvIOIQ3V+oROojEMRqnLOQeriumGynE3fINbTsTZvWP8pf42ri
Zd/5DnXy1mlp3T/lMR4UTVA2J5F24u7q03KOsefKdqQxEZkjz6D2o9Y+MLxv1GXu
t84a+sZL2wFDa1ACnGEO32CK+Ll1/3ec1WYjZgY7iEAbwaJ4KNm0szDYuMwGUQ7M
HYUzqkEjgvXo93b3kBlSW4Ejmw8HqStzHelHVg/jagtvKFFMVRK0HoAHxDRp7SW5
gJrwcp2SE1AvulquGtK64Kog4M2fPBWPEfj0KZvHLhiNniISQTRXbdzeOkABYfwp
+DgXf3KL6NcqbNlQIcRCNF2nqH6zG0nEglbSI1YakFBlsH0/JeXJwvrD+qIo0lBt
4vYqBX4BiMfMcvRZF7L59m2gaj2YO+Oak//5jS+iSbzJFlsBIY3tSN+12RV02wN0
tm9/T3kNep2nDYSWO4zSk0jntW5wy3OY5uW0ocVASw4mChzW57HUICQ77JRXUBg9
WN7A+U+sZJIlnjslMKrPgitLDetInDcqQU34cYHpuAMKvad0q04KdN71okuOXdfA
aVNKy9Vwb7IVc+riNCrbzKvTbC7hvgOmGStV9hb5X9Bc+hH9AHfjeJXakCCBT+xc
wMofrGm8oWZ/RvA3wsKr2Vr1q284td9Rodmcf7NFkIXfRYwo/PE+mWZjVwQUQTVY
EfzF+agMRJ8P3vMct7emIWg2rRpuQxQ5uZgzHLCa8vmrWD9gS18LruvRt+VGBWuj
Uq2uYftLEOL9+Y8P8SvN62SMRY0pDp6YA9XfcaEdU2Cjc4cFbpjb9X8r0IOlt+Dy
c+wOQ+9nLyGJV5SyGOxL2AZzZKGK10QZWDvgK1krv0ULFFtD8YSbHThr05PbL85f
OcoASL379oDuzDjctOPysoW/kgML+sNVRXy7N3Ye4k6jbLmKyFdb9/U+TDpvI1Io
2n0UL4ditVmp3oQeZm4XT3Gv3mUTpEM9hM7vXpAe1mvCzK1XX/0pV1sbWwpDMYP9
8zjLS7cbhhJzdjIZtKyps4rR3zV3E3xOI31NiJXa458nx1bQgYALtprb9nqphJfh
mceqHnydSQf/FAmHSvnwRZaIq/GnZ72ZrJWZePQ33wtwpkBtkyYFws0SiJv82R2w
NcJwFl9A1EOmqgHhQg6vyKP4Qg1rJFs7I1bwl0k1JI3yEKBM5QkewgK0j/7UB+sm
0Yy2tPBfCVis/xi1KmQD9MhBPWWpKeh1CpLKWK2CD8EZ9aiVgRTJOKWUDMWZtLQ5
HJq3lA9pk9xHxUscDRxKZlHbvR66NksRLEOV30BZpf6uQJBvH9pKe6thm4yEPuAi
DLf/2gBVHMvJ/CJPOQDdEaVDszPwBnREtFEnkvRdHtknPhrrQrd5PKTa+8AfxVif
hEktuTXhi+2+JnRZmlIMIh7V6DsMQMygDlaMhDJMSleWeTmd0m3ewewlLjzN6XTk
L2PC/0rghXOeePdCIPfANfHg2/yg8Whfcu3VjZ+mHx02MAYYeVGaTHAsygg9bFvw
DfbVdXEtQ3FDWIf2ieSd/uW+JpJbvLXhgBeicQoYfypfFRbaslQd3l8V7aL1eEsi
UjmAp3bLDkzeDmT3pJjoFyTpJFfTsnmcaC+j1HVEftt3Uj1fpZHkpxyk9W0JUcYi
4JT4kq3Re4nOMXyu7H81OFyG5yTUdnwEVMavYboBv1z1KSo2GFVgtPgp7R6p58aL
Vf37PhyC1pVEBI0KQXZR1P6wUs1pRc5xy/Bw4BNQdOkoC3pEJhVZ4aUJnf2a5Z7C
3zWpzSKPyS46Y+7wsMlfJ+PaGRAZMH0WpBaE2CifzVoqMStkWz0oWRMsDnBwdZd3
cQ+8B8pjKx41dR04V5VGYfinsJoM6IogZSfbW43AkwPyICaaAWO0AbnP1cWEIZJg
iGwpD/wqFvqp2F4EnSaA0XaypBC6ZC0WP9RqiMcvcmw0GojsjsE2NDZ69vi+zUIO
qU34hFWervNpjT802Z21UgabNvOc2a8aYFq+ewFi2p9g1WhO9g/PJmyXkUWK6zdR
ctepx4X8w0fdSmakisd1KhBcPWWKpMpacl4p7D2XBoIQWC6bu1QPvls6pZDvJN71
4945OjsQknkVPahoNVVSj1DwBeQ7U/zjO5b5mZq4mzUSIsoQFnhKALJBO4xpFOgb
nq5I/xNMGGgXA0BHajMZyxgI7vKS0wyjq+HhS54rmHMfzlydk8K2KKAZubOOQi1y
lfMvE6DDpPiLjurHxL16oTzFf3/8spK3btTf7SCFRWZUAZfzzg9NnF48qvVz3YAE
MEl9KEP1OJo08q7eb0VL/mx7bDKgZgKbP3y0iQREG8aeTvVFKL1Se43dUkFfU7pA
HzUkFq2NiUMHVy+FiEljSajm7JnfBTN+G7rSTNojJgxGNKn7Lur8Cn7ms1AKtV5T
bbU+HPO9Wl+uoIJvDYDFmvLr6Ww4OYCmKk7XzwtEL2XonpNFcANCPBAePOPTRA2P
tF/LlUhHZDvFarV5JoRRu9D26oH3KyjsXgY9pnp6uD+3O6gnnytofJb761tHU2ZR
8PoJnCDgwRM/1hOhrfQM7Yq5IRG9/YV5MUsM6sS+0jy6thBfVUN0Uv5IUImpwA87
sWLFBtwpEjwhrD/+ccdHV/RvpbOzrAhgeUs8plDTaPhnehP8rmp6x8TX5PL1ej3b
jj88T28BcG11qsHZH8kryq8vee3vZKcmxjQ4h9b0I6dHxtnrqMRe1sluef5HEROj
EXkxTGtCaeP0BjleBGlq28fs4Dg9qIl2bhF4apRgDgKuVTwlKh0cYxIWkhySblRg
19vwiGR7Kem4dWdk/cTZlz46PNvg9VP44/vM3qucgQpW6xUTtkXrfKdnn7tdrVaj
YxFKHBr3gVbG4gebTAKFnWLbRZylIEAfBYwQO+7m+RH1L8an3g59jSSC3W/F+zQo
sNnfIb6/rsibXzWY/yy6XmLvxPqEWfsb1/pI2Cyw7Gx2o18Li28NNpCriPewKJTf
pOwilVKakv3UzWsao1CCKs2yVSbSQ63h4mJKiUELTIlo3E2NRDYTc4qeOrOB0lEA
58HssCw7WSfhqiXJUWkbEyNuck/n3Cfyj7FHFWIYIolCNp1rYlBwxFbwub2ZsNHo
rEOFVDGCDnVCAaVUKTkhM5fhZ6FF6RRsGSd0arP/HncRWzm+wNvwb3O2+LK3U7Wa
IpFBPjT6wPkush6Rte637i8M1rDA3qwiG3osrSva33Q26glAfvLu3bxUNMDQJq3u
haXhcTEysh8btfGhg0ftW0vg2eGQs3YsazhnqOKxGDDcPs4X95eoDwAi3mLFre8M
eoD3kdQ87dglY4wJ3ZvRcTc3jlugaVlVAySDczf0n3W4fm4RoOvKNCtAkhajht/u
cnopOMX4mGOcQqZZf8IIVvJBOa0Rva3NtPjakJHikVZYjhNBItmK7yGElO+GRHL0
MK653wgAu/wXkdMd+IYNHKUs1BeOpGCq5/xNoftuaIHEWuc26VqolKQiPLc6CEOf
5LJI3rcZHnwAiYRNYivy35UkUrpJdSkKJavlZ09HKsy7QnlcdN5xJ3W4lz1HdRRg
Lli0Fct7Y0lL41h3NDL2fjrebRQJqzKEtTpF6KzRXamyybEBu+odtW137EeiaPF9
+zCxAKWQ8Vb/6/q9rgVjEBcxqA1lT+A4ZtZGLsfJJMH1ofj6qIhtSGcbaeTfqxtv
KD/xUE69wS+/183gNzfexHXFqHAkRBHgjKqIrpoY0Maf4etMAnPztrhgkbRwVDyw
Iqk29tDt7CZROZZ5Z1pqV2gCqcMKEjDB1Qxwc7/zzFKyuRnP7Ie54NGmwhQQB7Sk
08eoPc9bplYT7B/VkTWxb6VGJQwPgHpVlDurA7hOXudwtnFgHO3DZKkV7W42lHHT
g9Q4Yly4c6NKrUPD8QO9NYXzX2ALZFxZ/lw8+m4w1Fhk+gKCYVIKD5pIoorqBkfC
blNybOqMf/nuzVHHkjD1BmgAOkiZI/PibYoEmWKb678SVlY8cRVJ4tX1GL6kWA8/
l2IOlK+zWOR4BO/FNoTmELZ6EJI4S+QUZSC+ZZ86lBIG5nHWrNhl8bnkmirMNgB1
mLhBzq/aQiyg+X+kbhwnOnhgBT/YIdckEL0o3DaSE0epn8O3ECYmF8M5Uh2ebX9k
bv0Tx2viG16st9Ruip5PTydXsuLZidDJApkXP7nsZ6+OCxugli9v+AF8YUWiNbuN
TA2kBFCHN2Z7qo4USaW+Hn4kRbTSbVRUdr4bH1gFE8qjwh+j4IzfjTEoJvJgyklX
XMMbS/vjaSUXfoXHO3iN8VjiWXueiEILA9EeNgcJiOZmdBIwBl4gnu3xeXIVsas/
RrnWLapERU7HVgEkvgk88Cgv7vQeiZi4RVbmdddCh/efDsclhx5UWcVaznq5NJKA
v49q4nYEgTbxu9aJyI8s7uZtr1vI4W9Ikc4qb6qemZZTIWtpZeYk1KQ2gGIMhC9Z
DLgRjTq6ns46J7wInbf1bwXDxsoK+tiIIexZgmuedRI8/Wtc7RYWI9/k+GA0Ed+8
eOvL+V4lsJXKFrKGGXYwMIbLq13kUEStI31dhgt4hWHT2p8BhNDfGBLXDiufH7OI
Cb8zoxpsIyC6tpOA4m13PQ6nnrszMgeiqJXwmIqehvDyLKGddyQk2q8llWgNhYiz
3Asm9GquFrwX66NovIXyY1c68PxFgwSfGa1sM5zieDk3jSmvgxUdW1HA6s9AeXc/
ncfq8Uyf/SCr7/jCq0eg0fjn3XqK0AgfK1z7o/7WmnQB6836U2Zk8dmnSKvW9jSc
fAu3UIWKyRNlBl7wGqouwFzGPQAez4dp5jKfS6eC1UvXdsi+xToQucCxPr1udYBt
qO5plzzXpNBOLR3Jz+7ktTVwlqXv3YuweMhlxPkeyhYPpEUKQpzl0aUwHkqaif4J
pVASxtMExx2M+FlakpnS9Z6NJQ+FAen8pvyAqqPoZnnIPtg6Ar5XU0XNapv/DSDH
EEL2XsO2+KMHVYRZaIMyc89cCuJZHYpxRp+Y42CsQ+0jc0jN+oRy2XxG2BI4vgZI
RpcnyIZzsNdn7FfD+U/fZwKlfeo0wytIr1fL5YmkupnfKVqF70nLspYhvCk24HUr
386OWCaxqfTVKRZGpUA8rvZtxmJ75Q7C+AlxGcpKidGqxsjs1HUr8Npid07ETGn+
Wm52uZ+XNcDrAfay23kPidnEcWL47xaQ3y3xSIym3fiFDx+O2AW+VXAmIs/qfKgs
O71ktAkvGOgdo4iBK0i+4MCn6LtcLy40y3EzyQiEv1+xsVBZ/YRKCYiAsieD76SE
diaLhzUIEK9BhPzzpNpPNZcuqgYMSB09JuCjTL7UK6p7ylBNvg12/DE33OA96gjV
+oS7qe1I9KGbIlwpe/WhjKe67A0Pgz4ce6DPV6W12EDJQXTy4qjzeNRCPtw6KAsV
pmgGlWyN+rEjjyB/r57jGyYJjsvoABBdiTlxLk9eh+AIoCpkvWExWS4Xr1kojdWq
cdVGZjW92TAX8mDiXlJwabQJP24nhpPd3Q9hQxZ+yk51NvnPmD8S7vWT539+yD4E
EWYOH4G9tGI3swJwxM09LLvYKOzk4M7aF0s+mvzauV5cQLx6qWWMWg6XugeHAGrP
IcX1RmXnoSba4pPlewxWF1n2k8No2FosvDZB73IVsMxfknycqTSdvSihQGC1NFF4
xFGotoCbFL/hiSwr9asiq671omtuOHDBBQUZOme7LuA8105/7HQ1I6ClanouH99M
2PkyCIA6IGeBrPNeNK5oD4iK8JWRrNlqWPdXqPhpD6jZl46yEv7fU5fQ96zEZtUJ
+Psy7eJkrhH9+lLPcYVA1nvuRSOL4LziCJujzwwWkz+EkmNYw1tcgxg6ce5WnvW1
pydDSi4BbrKREhnVzyuoT/w7mH17BEashFrbXTV0BDmC/SZDLCUMZdF8cO0rD1uy
AAK7p8WLchRwK+Exw2wkLbFVGVpuadGQjWYAAVga3GTF32iLsKhSj5YtzPvCLvdl
O3GH2TdbOs4ZUBMnaCV3PiwoC2lr9loXWM+SxbRmhKUIsDbPzNKMN7dfyZGym80U
Bsv6xVoHwxgjuGOqFDg3YfJDAw+oexNSRg5XCI3QrGJDRschf1G8Lx2+oBFcTrMV
e1YGrGT0qAWm6MEmaGiOxTA3moZjDvAUPon5EUfijd1rVHWRKUzbNmMJNrwWjia9
o3fhsdk882MMnV1p1AGrD1VyY012NQSv7+FysiadZOANJhs/p5MzRPSFovFpZqAr
x+zOCexTwzjl+70U6XX7oy9w/TfDO6PISlQsvZ9Ac5f8i5hsSw5lIlqMwn0zu8Ip
CiD5fvgV2II0Dg9CcNg6ugcGROxFJCDO5SpU0dUjd8CUx0TqRZ1I0i+m1yQeczeo
5GUbW4q5onnShdE1aA5lVgeks13UQQQErNLDyif26mDdhIM6Ou8T4hpZu0V2M5gu
JjZHSMdm/dtGDQYqpPd1Fm6hGFjFfSs5l1/ch5gcb9nNbyinA/cU3g2Jj9d09deQ
4vkALRYyFq2OpvYzXmAo4/JhxBUY00U554xCyF7OT9A46FFg8qOzK74Ucufyt+Bq
HB2g+xDA2UDxVPRL5AGyoKBpBd+kWrU4BuP156qNoQkDi1UAyvo3Bt+cIcvn9UIX
AKXQrFAG10Jg6AB0TgUIWOSWfJi9GtJ/aB2oo2aVGuew33WZ2GKWaZ3ubMVaVNPn
Hzf19XhIdIKdF8qZtUSZOHTp8W7uc1lPu+0FSjtneEsMjIvSRNuw1IOJQZ2R/605
Ggpq/GB+a9PRFs9+VdH/Znsgw+PCYGaJgA4ITyFptQGTLR2HIylLIly+wWF7vQVC
YNnBkSOjVkF/3X61DEtqtmjtku3Kf/gMXomB+f+rg2Cf19RxTjUhGtjod27Rop8E
RTY1W6+807WqC8eWBOkq7MV0KR27JwAklrglc5JTFrxYmOW0dJsgeuctQgh4XMk2
qo0GKfBkHXMOHHKDvgRpWKFuniBYIGSogLU4t6jJsT7PhuMZMwB/xu4neCp3zPni
r2PJcjQZts4GMU7MkSoktXTXP+rwVcQn29UjZLbuSDJiqLrPlW299bRt014mJ5zO
EYx3miAYlKUVNUBmdBQSqVxAowDmvrm5jIHrXJfBTq2sIN62SJqmNRwP8l3f5bKx
u8CVK39ZeVD4pR8uPApGmrrDMKLCiS8wnbnbDJhAIYvXJjXvmyZ3dmrgKyQyHcrx
P3AiFIsweQ6G+1HCAXz1DCtveAzzYM2fQ58iGNthr8GVIX88gktmrNDVKwZjJPpP
15LuPvLgt8vH5EfHtqewYNm9r8CLh37/vAZsgvzDDtxOgHJ/eNlapF7gPneTlGC/
D9kW4LFo6bHDHskwEUbj1r2mA7kxhS1685kPqiGNgPJFWkHt+qTH4juXDfISlg96
NEIBZADH+/sE2d2kJw0ZrobQmB9yvypJ3wSmcUd/q8pUJTVftDdsTmcG4fLPnwLx
IhhXwIKuzLQa/doDw2h49EXVvgnFKCBhg8fqE6ECQyCeHLODIRyctlPWRWcECmyw
7Yb7s5nReF85+amitzUSsamIt915Of1d+r+Pb2agCRkOxiqupDhVSWZkhPQEaseP
78gbKc0ybSN+mXJfi7ca1yE4HTwVhHABgip+UTZyM9+GLqfEJ6LOhsve+BIWsB3G
+TDtqRI/rkgSXMT0g0MveL+WzkT1L40OV6qxGRgnXo69S+Jr9mv8hyJQtUwfP+Se
oGqaksMaDD1RET6C5eP7hBh0b26xmKOqkt5T/lQVMPmhvaUHa4WCXjybi67gh6pF
6tIvpMH86nVoqn2gKybnGKWGP2a1joCgKb44hHg7l0cdkz66WuPKvSK8de9ihTXH
cD7rRg1uT7sbVggzdY4suIEKV7kPVA3uU8tnxshvxe02uoyxd2td0Qx+lWTzIx+g
ZMwkXX7p4W0QLwJZki+VclpmRCnwAr41kwUoBar5imqeIK2ikdaSChhi1CFnkrsM
oOtWcd3uToiNFoINQk773R2WKNs/YXtmoizQFa6Pde8iohs9DDyYv/kF7mqbSzLz
MoU17V8HmINvhp7c8U9Uw+ByWn5w2kjIKXmYcrn3qX9ivAVdxcR6ao8SiQeNeRBj
bu8OWL2t78omlVdjL9ya0uwwAMfx565fmTeYhKz+I1j7R9omxGtHTKBPJ0JX6xjl
DZwnshRZvJ0eqcjjOfvIuo5RLT+sCfReqe2rhX292LNZfa+XQET36HYjeTT3I+bz
ekFfNI+INqocPNZh3zifRWC0dZITrhCkatw6dA2aNe7O3akznzauk1Cqh1wRHtS3
jTXApYxE+qocyxpRDUcy+iCMJHQcjjD/C7Bcr/q1D8gKipA3NypiQxs05t5q51O5
k+i5KRajBuJuZ/sklkwqX1BT8iF+0EErWi/9Faa+C7hg1flfru8cwbmB8DUBz0BU
Uu7WZM1bTeN+Bm7tTx9fDRnYSl/E+HuS0iGOxWHTA6NkrQTWXDdRpVWWscUFdR2i
KlMf1N2Es4uro9KZZ6m/8TGbI8xzE9Ukk553zT3yZRebSbUdp7M4iqOo7sQ6sl5l
CTdIXVU47O1eTV9cI8nwWdmc7MHZAqS7nUCZxd8uWmrc1tH1xJYlsm4sg6r8QGiT
5jaXRjshuurI3llItooxW2Jq3ym5+AdvScflPV9sYUslyITDqSQ04aHaHbJ7ufie
cotHVoSHMcHbTIHmh2Xrxefd2ugUEDMixQ3eToYY5kfC5mYBfwK57WAn1eE9c1na
moPQb9860BWflhKRqJ+//8iKpYn9lC5MJ0igcTEyflxstYw7U+QsMf+BqdZZW4Eo
yAc5yGCX4OfojCqlnM2VL8y6ymv+AaG4Zd10mD7rdtosoHbbxOgpzmgtbJz5kcVk
bOIP3NiUBRl60S1Kex4QEBOQpYZ05KSUI7XIlsiL7nrMGv26bqe4REoZns2+9mr4
496cGAVm0ClgD/ecdVwI0H1BsiOwgwH3vXv9wx/iGJ+BEZxD6iX/xKc0rfBi0W4m
NEZRx35I9J9UfToPHHMBKKsxhJBs+6IDkCJCsQ62YDuavN2L6Y4eKAyFVvZpW0Kj
t535ep7YS0qFgFRytv5z0WrbM3x2DMvM0FkHcg4USKyk3sV6CAo990G+E4QCPonY
hJDMlHL4kek6zev5AMlr81rOGEhApahfS+FVlpZZUzTyGys5xCbTh2aJLTun9ZNJ
qCvTIrqmXO5muTOckFpaIbwaoDmk6ErTcLz/nbp7XrDj+oB7ndYYWLTEE3hHX2Cw
0irOVtx+Ixi33CVWqANoZBjv4dmo7f0ThGYBrHLZeN7fgeFYbaYryUEKYSltIfyV
5P5Go3TfTZNjYuwJMNzq863F5tX1eYc/xX/ysGSQ1+R0gIPYALxWQUSc3Ot1mPQG
E+U7XOYM9I+CkAG+o2E4fwJUMR8fuDH/ONTmSUFKjgEw4qGcquMmyWUkiIrsWOWi
HzTT9EdK6wFa5+XwBF9s8CUi8xCpkD4AAARZJWOLyLaWzRBBhBb0FIT4iIhdNrfQ
pQuMBGydn8osAM0L+57fyNNXCi4U5kaxsS16exbh+b53Y4aeqS8QKVT06QeUazyM
ltrWpuv/UFYunTTBME1mhHTdGAaIwFnpxf+PpdwBQBtuIbLT1TYDwoClbKnwZWKi
5koggJKkYeLcxmQoL3yVmN4pNlzPyfLTBXYddryRcMZD+yWsbY/RJ4E4knZwZLUF
7N4q2KjfP8deOYaRd8bC7Bv6zAeL/tNkEfaKvxQuAPtmoDKjscwCRpxwdS/d5j4X
Xm7hdD3kLfMMetGIH69zcdYIqrJinC8yS2PM5CrwwnEQ970h8urUL48hdrstVz5e
RNReMJZeEZMwtGynxDZF17d5ZverZwL6xFd0NWt6XTDdy0h84bELH4UKQvq/A0x9
KHQSGCqzmXo3oMbEq5LsVgBUHfM98QMD0I3rtA0min8hzaPnPzoUzkF7A2q8+e2N
Z8VZ6az5QcQMRZ67sJKJpknVmpYSbLxyd94/MDJlhL8jnhTpFSkJN8Rg1ChBPKAt
l38JXsupfqgH3L3jOX6xowvDdbqbub6Y99fNpG6oEPAFYHt9DYgtaL/NgWwoB7Us
m3Dh7GgAAYIAx42VVzyx3eRxqVubxrdUvjeE067eq3BumgMYlwkOK8DIrM41sMBB
8ioqGexX1axoWi5fBHw/4CreniUwaEVcQ67RR/t+wxmhKPI1EuinX3dJoJp+cJ2Y
Hww6E4t9/Obd0gyeOZrERVX61mBWFHkTi3P6FkelKZshKR5Kj85N4DDPeeTPknYq
N4HJo/rQWTQJC3EGVW4ZvmTVD3VA9GFiwFqtyfD7DwDlYutRmzrIgPzgryh1PYnC
xpjctTqMc1WVimm5O8arTMdHJaRG5kIxnU0tXtsSa962zAanw4LXx/XSprZg74Fw
EEn0z6d4agr3uarvQtgzl49SfGbthQKbWgnYGUfmk9GCPAg4PELAuhO20Z/ArE3A
dPO4LsYjw/Rtxwn01DBYgtitydxEkAU+rcXUTg1VnNe/sQmjCvOFLKJpIbSaDHYm
JFTqYvBT0QYGOModAHdTkBgs7gUXRIAJxiw1L7r9Md7GwOFB+m8wwf7RpvqeTH90
0dUJt9a/f/S9qObkl+1o360ufoJPVrCwtLmUdY0vSKYKaPoUZd43vq1GegtWtM3L
rR9mo2Rl15tdEe/p4BfgHLBg1uRzxu9ZougnOBJJQL5F5je8iuCxhAIHsILgdp0y
ewzDNB7jorL4p7aqX4PeBbLTzAZK7+uHZRHYDueQ7Xd+sl1TYeJGIjxzHUa9wLfD
JVb/S8JuPk/LeZzyWMgnCX5EPZrvcOR+t98I8D4dnB9YeMakb0Gev3ezaMZa2ZWw
rBzdCurSyQNcQgKf4FCIZwo6YkswKlW5XNdf0gy4KcopoQlyloWRjzpDHB20jf7K
3+AcdruEq2gFj4J3W3AZtlOSn7N5k4GMfCQmmng1cH7705i4FiESBuJq0SosYZMQ
Qaqjn7AKjSC3UI5RX/c5WKEP/FcUkxnsZjdSCL/IwoOzSj4PnOz6cte6FoQemy/s
AvSSGumsWlRbcSr65WXi3o0AYxUwNx8MFN3RQuvz3UcKIGYxWsnkyFNfpxX2yco9
IhWhYGQEU6DFuhXOegJ6X5AMBf94F1LmonABKij7/nZXPCK+6pC2Ykganq+bprqC
zOyHX42nuO6ZBnWsxKIiH8iBMxa6sYJUCpBWBN7F0avwk4JV0YnS63RNtorfSAmo
nMnN7yUYuNPiagcy/GKP6GKdYcJ5Z7v60YKaX+6hqL8JaKQhvALhJB30uII+c6AL
b59UarW3a76/4Xv4rht7AJnUA8Sb3qde0cyFvpYyLpfADcWbLPL7sN2yQnD+K2E4
8rsVoFqMxIbOvJZ+T8OYFwyTTkgl3QiN3Bad1aZr4ay1pbIA53mh+8DILPJfPCaT
728L4qkjw/Yc/e6hTtsoFPFiNmbq0oPm6UXC5wo86lNcZLIAFyunRmfWPbu+SHp/
ezIzW1PbeCz3wvQdqjYx16RvxmA3suPlELgr5Hrx9bLVkvVuZvcrwo1K82HTARVv
+cmBG7PfXj+W1oC0jumfTJ08Jfg2JDDnS7/sAPsYxRgiUKr8zevPdEZs6QKmqH2E
geKM2PeqpgxfCtpxG4RbM9RyRwQhQIsbxNVzR2jlG8khWn9ldOCT2fP3drKDNxAI
bwq+PKpKEdGRj+3aE+O4Vuw8O+L2aWXqhZSN8Glo7SO+A+KE0Xi9LtJ0h14VpGiV
zzGDWiAQ/h7xrCP8cHtsdUOYbo2a/6Zruj5GqMfMwTDaYrjDk0xRrV8lMf8c3ml+
WJCJ0vg8XGalxNjY81CvQWU1XTgceMY3fKpnSMHGcX++mJZrH/qmlzcq3sgHLA03
a0Bkv5vQ7X7g08M6CdmekWHlsq+SSfwR0lK7cz+3sw76+0eZjrfpHZRHY5vDlhfJ
1pZk9IBWynt4X7hF9d9E3M8CMFqwhWaa/PcOngzMHEGMv78CwLZYuJPp+wGJIw2r
OIiujoaxO3Xhj+bcJTZbv4OTnGM57eyZEsUb8MkptP2y6cK5FNq1qx0QV6ocAhYs
sAiuwKMg/c1jpMYG2ET37tVIJJtVjT5jZqvk2zgyVks7byQ8OXK1qvV+16VFkse5
2jQhM/ZITFiDxl5a4zGwhmaVj+2tgnACDpLhYIXFXTm9UDusCEvd9KgOfDe67isG
fliwmwOYbB3RIfZYLkAOzHLYFH+AcMFmR1ZUQB7Yc9q3C969og7C+Wsw730wZwWv
nX3yLeBvrZj9wIhDfTiRTndTB4gdSJm5/A9yD9XtYSsTD2R48uykbgThwXXfDmYy
xCwv87ti/p93ZPEZoXjjBv5Yn76Vid/NiflZxR3XUJVI94YuRevF0KBA1OsLV1Ax
6k0a93QMGG+uq+s+YPl95TS8kqx/MtD/BxZzZGxjUzgzUzZfCPnHTuwks3SZy//y
jothVMFlTh+aA0H9VXLnjrgEbZhWtHqbNAPMkPp3AyG8XudimYvDPf91qIJwvW6v
BLOTCZtBmt8+tlLYJ18Z7IsVkr/CnsPsA12eife83x1qwzuZmythsqybOCbHolPf
QhlDrW+ir3x0gsmEMa9Na95yq+XJrcDNRR7kmxpTUzz2L7XVY5bJVunJCbttq1ud
oSRK31ZTpGfAQE4xFNGXSrxQpNkEgHVotd4CIriB0TKJ6LOhJ71vvsSQZiTLnYGr
qMRZ2NP69OPrxUBY6axY/1dQ4EufpV8ACGtV4cDOLRDoLYZQqXH62oVlayD8/Es3
r9BFgHeyamgznmMueOcNim9pquHUbj2xnYSaYEjLbOW0CaUcX9i6shMPWXpN0SLX
FP5mw3iaE7QVuzYuDMWRs3Ns2WiQ1CvGleuw8W7DVA53BG8OybOrBYAtLS1D1Y4i
4zGqlI1duej0Dp2KZE6t3DEdFPYCFJ84S5+en8EWiFh7vymuk52a3H8O+x5qP5CI
M4jlSpOYt1Oz/2MIMuNXOO+ApzCgzGFxiCTStimAjxwh8O8KUhBshtOQ4rtg+lyj
C1yJxp0ReUIDSOrwb2UXa6gr0+aLIVJG1H2MpjgzoB6vZ9+s+Pa50Fjcs+MgQT+N
q42hDuniYqEnFB8Vxj3xaOBHLyPszgBSelOoBrTV1caWp+LwT4zKfvtJ23yW1MqG
8vnGbqOe1aAx6shlCHv2/2gOGDy7IlkDDQHGkCWxR8e/auxE/t7E0ClP1qs14wQ4
m/aiBD83Zz/ZUNSgY48JEXBybaG7D3U8zz93p6CH+MEcCg/gT+VRLC+EG3DVOWmG
DQsr+e1xS0DNCxtms1Sn0TS3zpLqC6FCcISVKTKycD0AXZxI1/ZeTuVNzBQn1LN+
M9JrF048X3kCvInfXCjgi219yzMVKcylIrarjEEA7f1a3BNOGC5WyhNsQHA88cPJ
7K9QRvri2QRm9+60tCmk+IDWPjEfiuuG2VXoPMK8FhHnwjZTksFr8UNU98PIYNql
foVzHifQr6QC23acMnM32RJ/JQ7XxoJHPN51gWtPRayC6oAWUahQc7OxZKmRiLJu
CVgF69tqiIrEvwMwYLRVIpZpj41gdnJ/mQBiEaSl1Gf/FpoEuoQcNVYG7cGwaEsK
TtphdyJnVjsQCd3cXMx/7ZZuk23NmXcVkJndGLaG6N63TAU5u/mr5uvcgQhLvNO+
Mw1zImNkNYX2w6bcRRm5oenBdIl44jya0pIWtMGp0JwORqgmu/cxQoltoueU2JQ1
WQTIH7YjKJ9fRHf4QTQqVcv8XNj1PbBG8TCo4lk3JIaAFYNVbpF1bNE9FthokAqk
sQV9D99kcfVCfYDC9DjWDxk3B5yjmgrjqvxTxSJniGM014d/uacdclvpj/E68lXf
+bfJ/JjaPW/iu0pyQHgeXkVhgOPO1SAnsLOH8DIefGxCRRZkHNQ7Ev1VI1ukfoy6
WcrKmGhh1P8jmUlVqnqMby0gixg7Gz14Pk4ZprFzOhDZT+thv3h10JFyT+7bcRxV
W9ZB7Hrt11zu2GpK/1kacVP3UPcDgmXvZtu1ThjCNF7LbyE3jDU1E9yNk/JZYGtd
VNNjM3KPmmFAAdYx0x+c9pryivtt6ojbrskAACd5ycOMeXDPnd9uD5J/E6mnuUCX
toStJBaHluUk+OCSPqUVF3XqRW0t/ZgMRpOdaNHP1s73ZririGOVse7ToT2h4KOF
kNuON+tKfpdAx1ieffTd7lNHPoKOsjjLFNM1qbMhURzCeTvBM5Pgyk5eSouDfJQe
scSFn/Ea4CHC6vymTvtI5tM91dNVEFrYOUbAnPKhMJT7LsawjcJItPYsvZ9WZEuN
OTLS4oNXx8ZF3WAjNQTgyRPuNFOaC7LRlUz8Z1j2GfVeDFJAPowmgyz5osvOIHaD
eKwlh9OPlHZnDi6214wIgU1HhGZ6Y/KmW7uF/je14nRK5iunRXcunuCb5NDa6vpC
o55oVHCAyEzvByeJbiRc1c5ZBxqBK/+XOKSzxmGGhws9jMoF8eGoZgmE2s/SB6al
nnp6j54EBjDApXxvBHLEpHynZA/vxm8tWDtZ4CIosXa3FaMhMcSzkH/rA7hj+tTM
UD4QA4telkdekbbiOdYgnXFPRUwqY/rAi2fdNqS37bA/yQzFJlsGjBBiUpyzK0BQ
xsaV4FEh5ZlaYcnMhquywAJdoZn5/2nLryrgu1PFXBaJGb0tdcTqQ4ltLfzyUa1j
COZma3HdYI/RervlvAyfFpKeYu6hwFTYVN94yQivdhd9RgSk6Tc93ttoJmNLm7TA
S5z3aWDqtzdvoyUq8gdN2SRe/H5OY6rhf3i/7nOhVqcc+qgqhtjrK88//rebUEZC
+28M0OKpW9n+Fs/1KdnUBoO5lGsoYVzHpZxaj8R8VKx8tu0fXhmgccMg2eMOsUyv
Xod5AbsldXrCFow3gzCvjbEgvqJlvrPuQXrno5Pba4ahQUGIjSxdhlD5A0kqaDoF
fAVhk7PovYifuw42yiIhGbEFDtvqHvcy3UohjFty6jSp8zPdKjHObUUOZxwPefyh
hJwKBwEr/btTnzGYLdGLJQeFmo71n/hZjGZYqTSTwNjMc/tQj0Td3DuO8v3mYuKA
6+RLMYHpMBNMuAipFz4l6HTyTT0ZLBHOeqid3yI/C0lYtixzfhwyapzrO6NocpZM
kdrxFV306MVACj1Rn2m2GLXk8Wr2/SZpIA2EzYGQiaywXtgkhX6ZuBelJJmdm/IV
X6aS05SSpIqlVajwAZU9MhucaP4yHEbfHBLICi7oz3zYgb0UaSihcu2U32qUxEhI
7hTc70eYJP+8wJziZcGspevPFiAc6JUKS0dy0j9Y5MqOUaQ0cHv3B4wt79hIahO1
SfUaCHcF4/XUQ/RCpmQM5dJ60FnMJCMWovKFmkV/MVktPtpwOuq7/TN5GRqJqFMB
71YzVdVVGmuRgdfBZcg8euQaSlz10pRCQ8sZNinL5C1uJURjlvlh5T1xnrqyE0ft
nsdI3oW/Yyi3AzXxtkF9KXke/J0e4YKMfamtOkNXCCFbDOZunqUKcHfkp9YJ45CP
Pb4f0bypk7In5uB6X50XRCWk7hsw9XF4PgNycNeJofRPOTq5klVJazi3wTBzppmA
VF7jTGiRSSnHIp+dYtL+xsmcO+W9fdLrS21jlSED/8J+ofDWixZS9CNm9bOGmJ0v
mqATWmdqjj/Xvs6xGIJXEihKx/X7fppXDAFXbviEIn3aNqbZlndw6tw7RlYrCBRM
42UNe9+g/qkPOJxilPZAU3QvlB9mYzc5TU2Y1yOHnHf+vXYEv3v4XoskAF5jkvxx
xtapE0v82s7e4W8ItMlhlAghak0CKMrUXWDN/vWHg2pdwozx2zprZNSaG3LwstV2
bfX6un6jGLl9v1Umgz7ieE3V5ruVq7DzVrYCQZUrkAmbIOix6BlI5+KPlOnuRNIY
uq7RsiqRCP+Ufb86+yd0W1GTK8F9hNcZdrVtBsu7FnBPA/KHE3jVxLvjaB9YR3Ic
+tRGTIkkJZB/04CTPPxBFBlk6uxB4syg+HRaLjmLbvGfVcvoEoVLhIRf12lC9ki6
oY+jX6Hj6RZFMVfa/t9NzrmW9460DTgnoi6H/qBsK4LfADzMWBW1l8LnsS8H/De3
dzDKmb4iUc4gkabnRPSy6h3nJxAojZ4EyAdUBqyljLneBre8NKESqs4fjciycm/j
oxGl3SLomH1gFIUIxvxQ+jpSIuH9T+bT75BF1fM37rGKG9D4+znOKLtjjJk6D3k9
33Bw3v0m3uecE0//PFqVeCtqON+c9v+LBlcJ/TfHK90BbUH/swCcYsV2TNj70y7A
ZmSZmPkklPPtnrUD43mVzEnsYp4nPystqkNs5yIWHlw2uwqzrVQqssMWmime5EhW
/W8XKoBOnx4p7fEelgbeq+51qIfMdWKNKXfreTigwgKA9NTtEcb4rXgNd+/ICL5M
mW3wO+zBn/6gIlx2OI3gOQu1ysEiGyHRVo5zKWZ/JvmxsD5UblpowB0GOBFD0HII
wVpgvO328WhaXUCbSfqyVJFt8dQTum/Ber8FE/azNPXfP0sR+KcuGpRiRH+WAQJ+
bAaADNV6KFDwsGk3ypkODUuKvB22LXiEblDdYKGqnGcyC8WNoAPA++r7556EyEnY
C6e2Bg1juh654s8sEtarl2X09X3yJ8Wj6o1mtO3oTas7hiW4saxegswrpvwMxKvk
/V2+gkEVcA7bg9W8aJKcdBYogdOyzGh3DWCMIbHUgV4Ue2ibyq1JfVKeeF3WOtrZ
oZAw5V7hxn1FXLe0EDNPkl17B9ZXHqPoGb5/NgA8uH2sidIxB7do8TeSYGwaxmgY
//TzX60OcmOFYbzb0GDXQGew45TWts8i6wY5pv+yLoDYlAcYBEGXnTzt4fmxM1uw
R3DBnX1qdPksWvVofyM0oW4e10CHe7obVVSkiQL78KXXV4smodCmchkoajgyWDbq
0/yf4seAcsHz9Mm1OeEiGVUKnMB8mZdJPXyKNPVEsBVxCA3Ccnd+88kVvbNv6zsc
uVoeqqeui3yiMGNLk0ktRqZbR3bIUese3996ERaF8bePyTxgfaWZN8X9bC2qhbbM
k7pxQlBYayoLxJUls+QQV9pP026gUHu6gUP/H4Jdaeq6z6r024NdtSScLrdRPuws
yOpMKgiSBL4N9TQeUVl8KhFYxmb8qCY0StHVqAYH5yYjpQ0zMwN4w23rQsLzEhAV
1GiGPR6fjyLuhNVIeFrXIAv3Jl4mH9AMrcmbyEJfx7WzwhMVkKl3g4lk50nAUL6Q
X+l7QgtP5Hwe3JrBgEbkl2HEodC9t9xmjNGo5Kmcra8fons5NiqDndR79EdESKL7
/WSmQF8fcYsiotjeigB0suoikLs+V/4w2aop0u7jNSbXMsncFUb1heZZKkPDMkL7
7TaBhHDNIGDle6lPM1JDCrtl2OMr4txj+AbbqrofmqFQOBhDvJ9xQJQNtko9dLSt
A/crB3lntF2W5Hl5HEHqE7kdMe5ZxMPIzwI/dUQJzYfnSbH5190NdvgC3rop//SE
oU2dg12f9f48K9YqBfe4u+K/9UitnV1jJWt27ZPyybbCHYjEp+nvMreybUpumnkU
Ornpyp8ps8F0sOj/qG2p3LBqMoZZ358KJY8bch9SE15x/eu+gTcRhYr1UuDrdS/0
IKJNVMCfNT4I1n2+ZFaABfr788zPIobFRBuDBhrurkxsOKuNT7BuuI0H04I6czXI
QA5wNQA0eXInSEZYAiZGY56tjrhfqpSekS6kxHqXf4TE+t0WP1WtH837OnGGwS5x
WHPNWFrPdKcboLsUrNwinGGBV3XwSswrsf5NMC3cdOFqVMzqGKHD02NXPG3XgVoE
o9/oxtUPeOb+wpVB/Y7Z8hytqJB4NkSp35M8cT1Nf1xK0VebeECoJ6stPOglt0/S
nHraC7l3hnA2Jzdqu3aXVJVmJLjmAu7tTGlOuPCiEerGHvrlZ4Ri+dvX4GCDnAL0
ZwI9f2c7P6gXSZyjzvKItzih2WaSmrPrln2TtHjos7dOs4jea1kawbQkYObOjS6f
l7quRctvLPnoaKRBrAuWN307toTYZKsmXp7Yq/+ik6KEEIa7L9Y58gCJRWPc+BrE
TnVZq5qrVKqbqccOdahkzD9P0EgieZfIvp+afofUsUxx1rsinmPp7iieTS5LQXXg
FncaDNPrJyyKeEQNSpju1HJ2GmypmMsjEoibmEuofW4Tu22sVm7AkelTqxbshC+a
pPJgrrcGLCC8Yn78MzE/ga8vHMLxdAEYQgIkzCtKyPQj//t3CUqJWoRUhTwAglT9
WPt3ZJSFQyZJAIJC3G9l5vDytuG4qX3/nhMvnT17u8el69ZO8DqvUlOgYEi4Pcg7
rhQhbkYGmplN5CJSaoOd33oJ6qdamBoOT3SKvdV1CZjqr8+6WJimyk+BdKAnW5bq
iGZxGRx1YCrO5xVH0mvg2SQ0CSGDZxdPeEguS4wa8Et3ve/Q2LmJinzG7AFLqXdo
ZyCEGtIMSv11Bs6V3BF3sejfKGx2+GQq7aCJO/VcFXbbMqKSsi/AgRA2HVu83ssC
DNYEFFtzIOjBUFTVhI39JooLZFAVSLiPTsldRbMyyraZKLmQxmDcLLuVzGX0jTvt
RdKKGqKVhou0BBh19HYuncXt0mWg8ytEIm9fLWYotbbE27t3Yj4A5JK2yrAarvLr
uYWeC0A6QgHsW+gWcoyzjlu1Y/3DespzxVsk0wIyKT8cYlx70UmwDOCGFTwaPOWB
debsYUUNAbU6Q4f4jk/4Zq5ofXMniMNX4C5E2V89dmTT1Vqbz3il8wE7INcbYZ0a
J3yQUT87WhhIZHpwy2PNO2rolgEBwvVtNjv0Ed8NvYiRyAYTpqdC9WOylIlQLGua
SoHstcq1A0mDcVoqLsuggGU0DVZrAKEticdJm+VUxqSHPswtNvynhVazSqDO1E4V
CwcXqBeG1xwADADwuwfCoO/Gti9jLep65+RfE8X/4juxywblPKql1A0CwX7aFaU7
kXM4tUjduKSqYoOPruboBOZiGVkT31/2ugzZr6Z5EDGd8LUQtDYAqw1WzJ4enAGO
oyqaAfElEn1oPPTu2L7naF+EchgsbSJXS+klbkejoDGIMQSynO2XRUMz2FQXkpzW
x5bAYuHcD59QuXFOKQmpghDR1aB5+AS1p6/UaXgqbHURSOqF8oXcoFSsdz42ewVn
/C9VRS3RrGrFKG7XIFqFScRYouUMfwE3t9G3JUhl9ri+7v8rxFZAMiCjdVOuSJ39
DTxMqkwv4u1sJmCmuZVZRGzLHM9O0uWYX2PSXV5iwZxD+ha+LcyYSpT7EIA2UtG6
xsA7xaoOFWED5RX9PUUYxZVhYYUz4fBBgRDE0D07I7BzVDJkQhDuq2pj06PWz1IK
u1/7ZHNH1b9RwDkybolr79K1q0Pg0rmAgw+vaFvUhrI3DvXeDJrCxTmDPNW0N7pt
3qufRVa8475wRNZMa1cJTEpMFRfPO8LPA1cwVnXCJBRdmqH5FIy6IKI9kALWyxde
TLX49/vxQ2FFz0n5bsPHY/3Po3yr2X2vD+Bzv7+GDruMr+KMbNPu1aBjCIYwdRtk
vr94CBw66XHnOO0r8u/c1W6QvJOIlrUrBLfEl2bbr9LP8RVYZ2K7WWYsfIT5B78g
1wtR5AL8HE2RSwscTlzqmvtbz3d1S8Vv9Qt+5FLEgitndcieNIIg/qcJhBUhbLqU
sUuashB2t6ZRRDuZZtrJf1DmkmA8AU1I3r7AoezL0AVrAzvmnQzZZjktHAv1hS4u
/gwSUhcblDM3gG0ysEWBD8IYkkLs355R6/JXEQFJDzxA/SoWMzIfBF80rQX6jgVP
ts5wO9JtXa7XnLAyrosv36rIm5Z+t73FcpBhxnc28viosOMbb44CMGHI6C2LwjHB
iNXIJcHCwp/ECNEPQhIF6bGRulvniCuXjJU/WEZWcCnAOMc6vXpH6gFy2NBcVJXL
P3R9eIEAVrUTYIUMDc8EdYfnPSOXIOiILjiFZFSVRP2sMes4nmI++zXbbd9CojW2
P7sdWGwE/0gGw3AYxzpp6ZZZyw+tq5GNsOY54rH5s5dHdExj/cX4aL/BuKAukqN+
9xvfuaUzGQvLHbSMElQv3TrvRqaH+Z6rDU3VMUj8KDFmiFoQtUoMLpzh/SeOh6y1
l9vSMdSYRfFRVPLTo97UGWpJMvp2Wpv8v1+5MJjkkbLGKE69AB4ipYXu7XDY1EWP
4CPI0Wx0P4Hk2ukkGcbYKWT9e3e+QLEivB6m+oROVbsHGTtUi4bMQjfISVqadajb
Ei18H6AQaK2uKs3Sl0jF+oCC5+MmOpTaBD912AWsPGCZSTCyZqYegq6ce9/gtxAv
eDTdPzmKcMee1lfpks3VnyapQDq2bh5arCPPB+xSX683KSofkDdGyQ+isVImjil9
pA8Kj3G+Cah5w7rcyjgmLFMW0UQ2Hi4e0eVhUB3HzoeLjsWMmgyt6cvHnwF/lFTl
HAm5+xTPQ2exapiWhGprzknAoZIWqRmD593IUdcST7XloJWrepQ0A8k5M2M9KOqC
vlsy5BZW507FjipIbBxbf42g8W0QMVxLIzABaFXe8mrINxrhZyO8aIZvhqXcKRdI
AiNFL6jTaVd06vzVGyZ7vfamdX8mPe3BuVS098d/GdmtpQ3tAyadkDgJb/zgIrbH
yLOOoHvx1rGidNPrE9Kjr1ACHUznF9ou2WRqDemcDuCsz/x2UuzgIvIWfrHUqciF
pHFgnyaffPE7CStqafufSNmI2zRl6w1AB+8bAarui9gHTfR4yyzrzpaHeqwFxLsy
mYt5gjti//wDQVg+gr6Rg/CBf/h53NoxaedIEOmNmXDieDx1N86SjNdpwdU3MsMb
xUVUh7mkMoMZGvUSjmAXibFcLWs/HoScw4z26GJ8igov3lwYfripV900qMT/FjfN
tL2KZ/DkF5Kv5h7AoWUDFmjVzLkG4wG6fObFTP2z5+a14YaNQv4hn14EYV0/BCd/
+2fkncIyDXFjZh3cjFm21I4Hhb84zONvjwHrV1Lo/Bpd82BQ8ie2orYpYJS2mjmN
lQ8bKsKpFjl1C+X2MR49ScOjm1gkPhKTvWOKeOwONxLhQZ31cxHqbV8xytFXyCWg
PgrCAsiDzBzDGKV3+nA/kz8arlUlfhgu2m6wHnEaFErVguzSkzSHv7IygdYk1s8j
xLDVf+0/wE+v10aWFSqG3/jkNfvBLLhy7FuUP+fqcJc3aeNr0RyWJWKVjvtyZVJ0
gMBaKZMGzvbMhkkMh5yyy3NMmoU31pLjDiHAp7MwbcZ8eCXPzj91QpDpIJ6/Fj+V
Gn99me9HThuyMDywSNaCfpwA+BHr6Ef3p5o5SjvnXOw4guvmqERcG7DgHc85BF1g
w5EhJ6e/x5MBGd1AtplHVnjSAE/12GoxHVh2+XPX1hnXgQMWeblRTvdbsQBnOmdf
5y0FbZqCJvlFgVFqOCS1gRS8kPyLKsnVnbasZptGf51J8dYRqJInSJOAfty/VqWo
DiEI1OASmQYIRl3T489TDVpmh202iNadLy5t4nDvjfvTSMYpRLLqoHdhebZy8H2E
EuJ1SYylB2vfdROKgd9ezg62M/uS4rM7kApcuQ7pV/k4O3YzpnibLBu3LdxIQGAl
GCMi/b3tFv8GD5zdKmYJeEFpkR4Z9lgEVnetlQEnA6TS0KScwa2DauBIgfgarMi3
dZ/8QyuUNgK43dcy79XYnICUOLPLvHh1OJlgHr0OQp/2WRBLv4QKPyTxuIUgwH22
E4KNk+C46uKdAAN5kL3M215CdpfLgKoFYBq4MUOoWFrQdkGF6SJQCACt0V0LiCGN
77YbFOWbc79Flu61uyGla+SOYme4wuz39j9IPolgeE/OcJPzoqWfys94yhyxzKA8
wTsDo8P7NCjm1S+mtPMbfD/pXAq/Al7tpm2jD/Z2MHwuOD9CWLeltbw4xqZ9YrUm
ILPV8iUIvMFSV5srlWdHb/o2zUoV5FeNyMyn7qeewaEEbYKu0KbURYBUl3gTPw0U
2PU3WNKIVq9wQT+ksFb7MKN/dahiVAMv2Cy83Orrhmu12LidUO8npnakBxad8yMm
s4pkSS/MoCCpbfpnWprF2O9LfvJ5a4z98oF0hpfOrD08BEBFcX73BUmhUK8aeMXb
hA+O9CtjrLT+jvwidi/RQoMInyoHxQBz4/ngWbs83MeT9AHpQ3Q3nBBHLaYdh7P9
+adj5SBWQa8B6VO0ptpXOO1kcMIAoUcnH0uRUigW1HPeRFGUfwV8uRq7cCoLk3jz
oKbo/fyp4UIwB8Ok1O8J+Op9SibxhJGBYIhcNP7B/6wBkcDjd+b+/7wOYIuQ/PTD
8r/MbK8uEhWy7zCwE2yE3GrIS7CrN6qrL/5bDxxgzwMStZizQeJD49dnrKhPPrkT
yWN1k+eeGNErJsO+DATFgPIgGVAjCsZ+Yf8IuooEXEkMgbtSKw9BIsI8o9AuIljT
pBHJcQLNTqUTxX7dNVPJmhEKeuq/mKNCuF8BvHgt5cvjZ8llGfp/FOkMYuD0HF3q
4l+xzrbGxtjAVf4XAqNzndZoBOE2K3TonJyaJ+oAxZ6tfOIEMcDRXYYX+6viyi6V
bGPlDLp9gn/XAoUl3gOFiHnfWeXBFSIfugALglyvUD8RJ5hzReo/ENvPYTWinxyj
VL9vbqe5mxySlncKchQ5M0Rwcv0m9PNitMI95MTHNuO4guoJ1OKWIlOv9AeMkSCm
opp6UQ9d8IGGaCf5JJRGgwwQdUTs73Jjlm4OwROlXW5Mg5leKaNqZ0ZJYA9ABX/w
qMg011DE042F15i9gmJEKUU7JFQXYWP7fsZ6Iqq+D6JtpolLVvIveW6giFlyPA1/
9LtfwKpuHneNWSHtGFr/CeQ+BAJm30teaqQq/z5ipQIjewq4TOLdDo9LaR142SJk
1pW+mKl8xnbiAzS6bnpSew7rbD03oKn+WxbVj6GK8hqxLzA3ZtCkTcT9Nqujlsy7
np7HEqVieQJdCP2dZTsi7+j0SGtbEhvC43cJvrxgbSXDBwX50QCjXwvOPAX8Izxj
yCfSc8hRGblrdIHa8nAQeGL1uiqlx2XbfDS2Rah8/z5QGXhVQmU7dPgsRq3Jzl54
A1ICpS8M0PzodZRTUxqeNoNwtOBT/Zd/2NmPKNHvQIWtJqbyAyk3pTbrfiqtzCNX
WaIh9AYpHW4Craucbi3L//djr6mBVq2zyPQM+GSkMzZWzksA483p6jgOFvddBA+y
znKzcbJKD0WrDwNVImiIQ/KAWXmdHEgiwHbo2Ad5qnh5oi4sOFp+bWlimAuEsxhF
ymaPO04x0ib5acxBdgn1u5cICpY8ezkwxrsMatY9UGbXFacjoI4lBnEpCuOBmfck
jQPB+sk6UeRBIWI/gSKev3Ifxv6zYvDEZ4uMkBqb73gYZbe3IDWJkcoZHoaS267s
zehjaTB6XgXVH483D3w/4Kyz3kD8ik+nXRgl1FqPw71pLEuw7cNodQGdv7kRmFRb
+mszdQdHgSk4i3t7RctIdFtnfM5W7fXlQRHd7wE0iggKtBY6+hrFLgm2XajpvWGA
/pcsWeYMPi7zwffQFXO4++6lddj1Sz84abBnw5/w49maXYKYmjKTsSbAYU6e5C4x
oym3zfNjHSKC3IHf/0KScCxgza1R09KpZHvjwB6kESbMtF7NTfSUEpP4vlImGoDp
e0YurTERNl3I9TjhoPPNmxOG0IaF+zMrLZJFnote1aZo7YbsRfQzw5ul/TOJHRzw
CP22l+jZA6KErWM34tkaDC9rw1gqCToc8/p8jMaJGJRH+gnbGCmQ3UmUjLZPyOVL
bPB4wRr9a4RwtyaL5WCHS2OrZ0xLbsLhySL5XkFv5VL4Wd2yflz/h3fx2so3Woam
HMS5CLmyXBKCpKwsweiJ/nHheO4tppiHGWZSGsp3njHsSiixmKB8lBQTPaLPeptp
fBSe0The4tnxoMneAgn6fq+qCB4z+gHIFc2/ayB9XvQKTnET5DLiRwKhFUDSZDSc
m0E5A8VYIKKIJ2zqH7ikO2XS1dXnAW+lu6j4UZXBtc+ot0ICZiaea/lAiPB/XbG4
JFJjca3D7in+HJUSfl+ZIxCsMJv8tCgtM8lqD/UFVn9dJqojFWsZfwjSV1XTWfWI
q+JkWc7mpake4XDuS5JUpqYsI1ovdFc737Gu6HJv0L661jIVubgkgkmFG1L+NtST
QnQoRKzeH49FQhznMrAHJjslAvywfWFFz52gCwQ8kunIrSVSebN94udeUJhtjh72
zry3mhOb7VDxmOtnq/YoYslN78BUVJj2fA+BXYMTxePQqAmonenpPOnyWUuajJRG
3HenwrOv28sjlnyqwJPYPqOb+INa6eGk48Mmet35katpJZ7ifhMKVJubhs82tBQM
h+FWwiQmHGiZdR+i9dCArp884Q7J9vYijGj2amUHG+Uny1MO+B7VX90geEaRXMGi
Qh+wbJH9y74fIC+rLIlck/g35y7BYwVlDQGR6ZfTddNslYGm1851wyYlOi3tP6ll
H2PPD53YKUfpbzEFSS3dR1luahEWT5ih50B1DQlX3n1LU6yZeryZKy1kX+fRzLNd
oOdE0ezNgLGESWlUXsWhxrQpm2ox6mnyyNY1FZik7f+cbfKCcg38C5BCBIA45l/w
AlZHOk1Qchb2SuRIAu53Gxs/fA5L+FCdkAriCgy7qgMeJep0po4SGWdSkb5GscK/
wTrTVvgTkJ6Rz6JAsrWekF9t5/QWUeb9v/A4bx+irYqFllvzEJMkPMuTyU3GiemH
b3PmueKgl2hL7WYF3djAh9n6WNV2a00cA4YvuTxhJ+H5IFOGJcL8JRyCfTTVdKVO
ViqK8lJM5pebB1pfmYYFHpjmbqnkqsbx32dXpzMe0BSAqQKzzfo+7bS2462nc0cD
PO/gmyKAgKOXZauMMBiZrcpQKFD995Q8dt33tDGl4sc2H4P3/pXTSUxB4K624t1w
DjiBUMXsx9AYuJUFpWyN+eafmJBTOVIPyQ0kKuNYm3kT8BP2ttfOVwH9fd8qZa2P
9Cd9pNe40QNzOcPEgvkctJLF6nwy7ztMZXnkrm/ZEXh37fo+HON3ycK09Yd972ku
aMTAsVP7TiHBAsUslESVkTOgOjDR4bTsASYimeuqRRpMLXYknEwQ/TJK1mR/OvXe
L1c8H75CqEozmh2TQsL/8sGStWKjqo6+SpHLdVW8peay1/PceDaf/xCjRjTIa3E4
hEzm1aoi4UUTjMZEkfiFgfNMDrukFGpUKf2xehYHTcuaaQGENLGfI4YXxIDqI7ol
ykWIVZm7q7TbxvZOg/dW1Mff/Dsc4Ny3bGVbiczckuJ+K0bRk2ZY7nR931Rh4gYI
iRwqI9B2HUjqiXlIWWi/3RYHThUZE9qvJtiP6FCeIn6V3DdIR0/udSyF5UI6LbKP
TroOtiT/PMfXPwkdEJH1w6kmCFxuyJonvYnu6pwV1WTpwkZtyhzyp0Fctvt7YyY3
g5ID9oSNZgbmOtDoqNhhQ75mMBhHjm1Ro6HVAfQPoWsDe6NYHZ2msHjf+hWF65oQ
wqgoJRBNvT3bcM4O6pmc3a4tXeUwymW66Aala1x35HyRusV3oaDl0EkDgX1H9MKS
1cJQlUJPE4WMAa8RdwHfRAQnwjb+ESaQ9OCyVLVCXz4uG9LXtosxafYZDaRGfePu
FcQiazYENRpwM7BjXAXaKqI2pLoe0VIgsU03PlZJjgfoeI4qeXXQlnldBlZ0kbMq
qJCvzJAhwVFo2YYPtugemCNJpwjKvqFY3OeEbBq+I9AYFyTIenefZcTbCpZ3IFGe
EwjMO6LIVEK2ttRydKb8MRQGuER9LYdzlp+7hfsZn7XjN5DSSPDcK5IFI0VoEmQ3
kRXYzP5/veZ8OwlmUwYw2VHimPGc2NHv/AoRwL+GOpafSLoIl6beSPFGDru0cvAS
VgCDn8SPdQGDecMo20SbHoGjfQDs8z+89o1A0JN9RBp9IuOxSZpBvkf2jLbqU9K9
kA6PKTE423kEOkWmkUFdklZcJGVaTT8aaJkZBlo0rp1jhEskqM+G6PT5kdCqerBU
7QcYgx/54ORuls8sKwHcFYPGFVLmj+Lv1me8AXa98uC95OGp539XItobq3+EF9r3
jRy2ozbHdCxqIFK27VOv6ARP+3G6CnB6HXsqIBXY8CuUNN4o8IfeN0cUQzEQNYyh
y4U2Q99USUewa2ZoDlFdpZTyv7tSIkA/mxuG0Hlq4NA2spaPGj2WKiOLa9o89+ww
gKfErOlEpLM3yA3B1g5WKRgKn+EDrZhjTzU8douCEtmTQTLsLM3f0M7PZIh/fGuv
Tg6NtzR0eg1vKHjgfW/Qff/QEycLCHLM/9rU+syp4Ew2BZ2t1JyEFVAPHxJtCZs9
MRDDx0gXAbDowc0Y7g/RzAzoxcSftoB6OGGJ10KXd3yIOC1eZR3saJ58Gu+Vd3Xa
Rsi/uSmpD/+VMgxyljiH6Io0ZdskoaVTtOVQa8OpplIWS/78/gIMlQ54NGeRiQ3o
3x/ewAgRglnZwaJfuB4PsNalJSroPYLQtay8y6ycvaRXetKQxAguPLoCaVr8rnyw
musBFoLU54IG05TqxLQnKE90SiBApxWzXjbkjBHG9/C5cFUoMb/3z+28TO2VG0xK
QWTrW6aMvfjzKlB771LRTjl1iJ56QF68l4VD1zC9r8fkmA2uiqEplu9SeMNFoNmh
5s1vlG3VnnoYbMsnXjespX/ku3zsYfE2IEBhHprhEGP3YNYVYICeXNkp5qIGQ7oH
T4bFPY81oB3D1qcmET21EnBA54rstCyBFcaJKaz/m13WHrfcrTRu3AJ+oTKhVGRB
RafDmY/TYpddTW2Il+O/OhHkXyiKMCoAHtVdmGDRMrQIXZuVm3Rvo9MLR1L1T9MN
IrAZ7kbqkKnMoalaM9L4tRFKMMcP2S5C5opE8AgrWvDLWAh/TTVtBPFlgx8IUVGW
gi/+qdlyzSHfvlUbOUIMc1GOkMlUQ6XvxWlW9mlFN3mN48X7SaqGeZKJLbt/M+fZ
dBhGeL22WJfXkv8w7lR3zotLb1lccgw3SGKiWrLqJXJk0St7Xpckb6xyorK3CX3P
Z6KNbxk2T04PWsy6bnuEJP2QyRXLzefWBeIpKO/sZyGvUE0jzdQlLnkudC9KA/L9
ynXb2H2fAmdNV+2vHJwVt6+cwxcWlQBlyx8f9Ltc6Gyq+0Zu1fmaWAaBBIcmjXwX
4tP1ZOq18PHGgWn4SpFGGj/WHGSqCHPi1YS+aMrAdT3hJBFXWbraX3V14LgTcBeP
GEHt8JB/aCRBgZexeGaL4v/SJZ/L4LBYTMszMm/hZktBO/28KAg4glr2iVZSSB8Y
63LIxHtzs6G+NRw7wzXXYvfDmgR6MToAyTbBBlmMwEMIeWCKcSvXObJKlQ6oVZXr
Car62btIn791+IpaxsdXE8M6CooZkFxag11hP0bRkn2Ceu9f2r9/lVtESQc2eA/e
3vDA8G/aYJDKuBAFcqB/nEo1O03tHHYvve2F5A9KE1ZWKjL/IAkBSYVyeKVuiXmc
fD69aMEKPICCcYXmstSBjQLr0pY7NYG4e9B4XYvt0+ROequfs2U+7VtmW2jgvXXj
V1RTo/fqO/Aul9zp0oblnJqZyK0CaPOSW1C+KnXDhlT03sBqs3QKUYIbBkGx8cid
3oJ4qax56e41AvkYl/W+RATogJZrt1WHODmWahLly7mh/grPPQqXx664RBM1sXkM
eV+4WAcTBX5Bt3Byl+IEuUnQFW4VRs6dBpoKKnIcJLesHSfkLG3HteYFQap8E70w
UUwoG46GyRNFF0/fIvzs2865exGtFCqMJfVWk2FqdJaoAobfQhBuWC79+ZRR3TdV
jugtpXACr5rMIwmV5/6i0PbksxgazA/wUUN6nXCafmlvPSU+DRrIptGigi2fBDkA
pXWnte86Zmu1O6lFCXbphWAm18R8vBiRwM+dTBtPmFSMVzdiS6UFleAUvOZNC/fu
aIoKn5JBAdwobDj/QcflsSZCLS5xA0PDddQd7RapG9QGYsW/PsXC6eZ4Z8iDbCwn
jxvynUWgtpvre7hOxs7fhnOT/rZcu7oHoOZ60csjCzpLk03wEC/uqj4c6He+GQkx
5FzQ895dFKFGp25ThAl+Yt0MUN24r4QeZMIM9zex7+vYbKryNZiY93aBhoKjqZoG
OarWd5HoFdzl1z/PR01soJQS4r/vFaUdI0+APcMB/8j58eUE0fKGUQX+8zCkIBlM
j/wWfeQ5g388TOjOc+JOzHnTDWAhvlqufzJqRrwczysfN0khdOfbwP7lhNoXPm64
r1oR5S8CUp+jwhVBP3S8c3as5a2JcahVHw0oneZAY/J1gherNgy5QtezoRLGmZLb
9LtVxd19FjoOXjaQD1opDlP4W7w9XPGQTu2SAc9PYxHPLBuXFPKCTEbdAr2XbBKo
l790a6ApUtqoG9PvaroRHQ8X5dtUHDay5w9Q1UofmJLoXv3GTXqCwP8xGM9FYoqR
aZ4NkPKgHf9XbIc+F7m9VRYyMtpRCQTMb45lSY1WndQ8qDoMntVvL2iwuXnPL2vl
GsdjblQLkOml3pAZcUFGclxNFkDxG8Yqe8pUE7cl+saZ17NShwXA23D9qBdMWJt7
PR+qbtY2H0+3dBtChvoC2L4/bqRYa4RVgRaCkgL2noXqyEfP6MPQJlvP15emiyvB
vzEuTVA4lwGZ9HDbDoWORaM+WihWnrPlYPS+InTrOz2z6XtACvpjHOJA0HxaqVZw
pFLsdst5r1U8MvS6soJKNv64tS8AwVlLeBDe6yUeRnWdjmgX4NQQQ6lR67Xeq4kj
3LNYNYZ/kSeLQakzNo67/IBt5OJT2qlHccO6WQzWEAbQXNgWXHQ30nhgT9LzO+Om
1g095UMMhV2AGP8prPsgKBRCzIUMnK0IUt8D+x/0pbogNY1Qv4XRFdDtw6YB1fBJ
e2aIHzl+kClNouopnRogUoQ10clCyMq9MWKs54Tb8Gwj5s9BIcfWyAoMI7vobxHY
MgsuSW5iVSriqoJmftPjhG8Am61ZCh6RnpGZ8W+bzaykNb3j6OOdPXlMLMe239CQ
OlYj4TzlE2kSbRtG1VslIDqezojlHvIHx+qez0PYlLHbpHGyKqSJnqwBR9QZnvgb
PV7QwKTXTVfnX1+TCI25LwzgiIOxA8sLoUQZX1TVyq4jK9OFqQbL/fqnmvawuyVs
xZVAok+JGIpHquVsom2Dr2sKLU8BfAX0Ec+K9X518NKiOUe2ZrKrBV8fkZ1AwL6W
g4uzWsSnee6wmjgEexZCwC8hTfzp38TvfMvJdd2ZepsW5KaXnO7a7t/yRxCmyMId
5zAPBQZp3MHeORomkz3y7qptYgWQU7NETuy+RZjbO397OVZ5OM3XZikfei4YTFHT
h+CZct13TrMlfbsofH6SuHNxc7fcSlIkpwCVu+5m4sWRn6peCGhvmVER4zZLZFf1
rnVZKq6kC7qxNGB8PAJS0o+JZlQTKJL4kojUbygl8PIDZU8PFovs//6qTrpuzuaP
K/gIcmAoRyf1gr6gQawRWeYXh4uUkbI9mf+h3sEpT+TDIuVCJCMIjn/Ig8j/WJSU
HHf6ZgUSAUuCmVFUicmU31E4KAr0HxVZ6zmSNY5lQYERQfb7pNfQIrlwUimk8e6R
V5w5h8HmRZZ9HdFSCfmEVX+eDXRjqKox6goArn9a4/i2Vo3I2E5l8pkkRumBnZC8
HhVbaZMXgnk9zl3YqlBWotGUA2Nt3gZQ8Ul3fm+4k7MAHbpH3jmXx6sx5J02++XR
W8wS+IR81O4p7DFhgChSbfcZRhUHeTuuNPsp0uB1dxBiY+TFQi88lotIvrSFtP6O
ok6ySTVRdDR0/+8cuLc5UAy97PjSH9WRK5eC1ImgcRypuxNSRLYeBznQI4jdOgWY
mOC87MGXE/cF73CHXCjJP0bOkIje/LzI9U2n3Xph04/2auRXFcuwIttI5I66GZV9
o/nHuiPV8b6+3u+c/k5K8onuWgC0300eV3/fT3GElB+sFqZCqdb/MeAn6j2SnuWi
K5cvMjYWrdKfNvZteaOkrdMcApl1NCraRls66IbbrPAc4+f5PPvmWWbdXFs5FHKD
Rquyba/gtRG7ej6fZrBBf6w13VxgTp5tD6/pki/JdYCJit6iVVm/BGyUmM1Tu368
7gJbPOsURRbRrlmUpqmP0RNhTYhxqBcBMGYiosE67PVbb931tSfvAKUpwU1vUmk5
4p144rCwM3k0C/IPyIXR6a2miZQFxt53HobdJUYHJBIYDBcmo2NmvUVTwGnD0ske
z3xxCDq40GMlUMCGP4Mq/PCEq+Fil3nn1aIybynhwaRJfcRVLGWa5xQSIaVw7QwA
Z7hgsB2Lv4sINjcu9Z0bMlSH7hC4WvUSqLM+GvNxge0i+1b9hi88BEi7EBBFb7iJ
KT33UIh75Feu+XahUGM+c92PWMrRZPtemYuRe0Co5cZzXgMh3QlfVv3wTxBkDi+v
+0P3Gctn25zV0JVqhhKHgc4l0+3RzTXoLH7oaECGOSU5InKoARDtSx/wDdlwJpbf
2qnR6KObegL+9lxsjkwskCkkoA6n8wJq8bkTz826hxRywcaMEnZATY4EkJGnlg/W
WJHvN4KXLZMP6P9jteI6fIqX1eikMqjlb4879o2q8wWEwBjpQ0oaS3A6OLl51yXD
kwHyk7HxjvtI8c5M1FKsgNJKnzt0VShtvW0xHKVLiRzQ/rAYuenIJChnmjLeLPBP
QyFddOQ4NHy5ksvsRjjBoQcVvicK8l2yw6LA1dYHi/SmfaoTDkJpa7bNROB0pCBj
Pmu1G+NlkwJe0LfDbNBxrteAVgnDHR3NUp8JOu9F115GrtmfbRGJgxn09ErK6xST
R6IDNzfMWDw+PbG+NOxPYAsmagCnagXRCYJT8FkeyBVnf0h++5MYafrAZo5Do5wt
LWPm92f8WJm/p8uLYdw48UW1dWUGiosTAS3tYFx+fgZQ2wj41yENdVcHotLTUBlF
XJPICt6D8ae8bR/m9P6aPnH0uO4Nsi/8taODNjmzs3G4RSCbEEB8rOTjGK4UDff+
ytqitE7jmIHl5C4ydB170hmruIjOxV7L6/V8GcQpg+FUzJ8rncAn+QkfI44nc6b6
Q2FXj9ZMOajYFLGvaZ01NcDflpW4172CKiHt5QJPSb/zIGhfzCczZMP/RSo5kpNX
5BlOpwL7gUQsaw7Uk8csI8L9gW+Q6ttFPqDksN7FmWroP1qf+3OncCjz4F5CL3h+
etXNAP/053KEOEoFAJdmwshvN1HT29x0tbukJ7d4G++VPrkuzDXn1yZ6tsa8tnDv
Y2JmP6uDwG3oZNsq+HGFXTzjgKN9uj5+3HvY5fJ/CiUVfR96FfaHrwXai2PGgH+1
wdcfOa4sPayh1lMIiBe4LV1V1IFWeOJrBnitXay82tuVij6nlkRQop4MpbYzWEj1
llA/HAJkLm3exQ/UhNnG6MpjC5Sy4A1SDQBUjhWbsamPEgco/peEOqShAXddfHda
2Z/Gr9lBlxNQINGbexvU6x+goNYRrsCBlYy7Uw4nUCS2+c4Cay8+3gu+EBSluGFk
NS22WtXLSe23UOTwpbae2wqxt4rK3hFgCs9dzMk2pBQk/C6GzcnDVRSjD9XYsvBr
nSFSLRF2iV0NvXzJ59qwlCZwqWeVi94/wyZEaAZSNV8uih78G0gQy5BxnUFAAwVG
kq4WvVQ4as7v8nfZY5CfcsOYP2YnPe0efO8VoBR9J5ztANF839V2DIwZG7IrlvcB
B1fCw18VUO9cu+5oHaO4zrb3bfWMZN5NO2jBeo/V0R8KBd9D2x8bJ5U7UGnN9srd
mMgF9TfNP/N59z5jZUHFUP4BYFuSZBPE3b8P1i6V4EjlBXWmvmKjy+i4P5mQl9Bf
py9gOZjjAASZnwChxcFbquz8IeW7K8XM93tSiXycM6Zh2LhpWC6EskNXWQQfIdXe
YozUJ3r93lbCtdD4C1W5G/zyArm888+0h/jF0xKESqL07YvOH5dcCJrMN7IAoZt3
Ef/6MfGGkU0GGwTJxLosfvjMq7GX1U4zvZhrJ5mw36CwISgZa1PPY/ETwgFS5dYT
dALUUb20QUm6oT7HUVROivm10Q32vMBgVnuoJauj4nEd5EGmk0FDuK5CxWhULeBD
9RVP/nVZVsYSu6+a2PNfn2y7o/9qNdAkgJuRCHLe1T4UmJt752rfqXnvjcZw2vPE
vJCRk5AI2eO0RtNTIo5yqekNiHQikjZweCvHQKFfI0oZ+LrgTOQhWH3I+wpPeTIC
fP+YRGUbQxphZANU5rVDDBokF3Ka/MMYOVyzT/29ey3CzAzL3Xrf1NZypNGqc7RO
CziWrFg8igcVGrCO4mEQlYybDAkMRPkjieTRxzMTmGHFPkByXpAg8vJNw96a1Gd1
baRDplqzy6g4ciE3s2oZcSQFY75/LUeuojnjs1VSmXgXnQROS0A7vfVRsI1aQhEN
gX+u9IoTxiU0WOdwDueb9VHidL8DQt/Dh2ljFyACk+5SiFGL9+RawcGwYFpq0/Hg
CeMTmC/vo/H5dP1dPKU6y0bswskR+rmo/GMbPamc0l/kJTcM8W5f67eGaDUTr6S1
UwmLB5FO3XJ3y62EcTKdmflBIszaWDyOvEGT5JkYuoFiqkhgBfPAngbYSSQQB5S5
RaXlQXm0tB9rXb4R2cJSxdZOXzGHdtu+AI+yj0Dd/8AWGQUNYh7kV5Uug00XIKPK
6Fu7jRWhO/AQup+DLZ4re3PAvv0Ip2Wok7em8qGIG1rtSLCEzMo6GoRMUymth7UD
1gZB+JsWSVm947uLIM0YyaYvqkwCLXR1+qHeKdAwH7g55J2sOmpgvu9m0Hcxk2r3
z02ZSZG6L2EFMoNvgmUMzFVEFXTB0EVLTFkJGxtM9d+IbqbCRdNqrlu3uJBmv5Yx
IGV1oH9wdyQY4ZfkJURPVx+N9CEJ3vH4oPuAOo7q20H3Bmc9vdUggXvoE3n0/QPE
L46VV+gVKxR8/yeMLXpxU0Rnz045V5iYZzAKN/dWZVga6nvR6qMEnbKx+VLlCS7z
gvOXmJjeIl5El8CFwsJavBhh+CJ7mcl2UB5T3nnlSO+c8MPuNQMr2MmbN92rYaFb
eiiYvqdIWbXx9EHAtOSSh2N/kpH921fZb0OKwD7CRUZtQd8iZrGG3c2cRyHZXa13
Zc88BtSkywkOpYZ2eIjowpHzqqMLqWW5aJXXOADXlQlwDS/fGUJ0vE5e8dcXQG1/
Gxom3k/OOzxQNUAjqkn6vnyF9cG9ybOtouU/OjlZT0OakcwbxV/1XwIT1THNsIOT
F+zw2N74/ag6/DcXJyBgRHeK3pXqOgKXgA9hhj8Fni2Rg+cKFCE4o198mLSxVnlK
URGiC0s8iELKNQkb9JWl+KXLF2OAErfSX2r7Cx7NYOGl26BdeN//xLXuVcJf7kfj
zIX+2muGYW1Oc3RqMJKNVQGBR3WaQGEdTazLBWwEDhgT1KJ04vsXGLROA8Pe15HN
NWf03YuikIF3JMxFy7TFJrhrR6sUY04QvtJgWa3Q9JHmYvYWnCImjhQ/qY/kxfgF
VaMbEY+8Cj6C4YVhcvjzUsn058Vl1YqDZBI+VlURmzk3XrlT8tJOfGRxtUk0TEv2
6wHpudIof9F+znvkjSZjHpeX3QKwKaAO0b5iX+X4xdnGAvziBGNacnoJzg6c/ynv
ZIvUJDnwz4yWxrnmOwaokT6vVYAs5ush7FSDhwZnS6ZEZCGUvDBaaeuNG5qLL/85
u9sAjirc3IXc9mEsFAcTEg==
`pragma protect end_protected
