// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:36 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XQ8RBWiyZxTG4GzLW//6GpSOPsxY1KG8oCB0qSj52+UCOOycDIs6iCXIcFTrh5T+
GFotj2h47BHe/oPC2MjLUEUviHwPlsq1NfUUckxZOCuwBGWZMkennhQKuegjHM2l
lx84NiMHdFW0Z8LEaQTAK7ZUoGs/r1JviKNJepASg0o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
AhIldtK3uWta4qU6j2tpolDuAx3+ksWPHdCVeVqf8Onhfly84wSvG4JafEsNY14N
z+oG14u+lKR4AdIXuPDrocI/+OhI3enOboSMXCIGeUnZ5oxKcC5YERxzMUiPvpIX
vydq+Jrf2U+s9u4JbxI0w12DKlVaIbFnKzWp4u+qsTjtmPtochj3oGWkB7Iyf+86
d3Ev+aDzls3lThjf01khcsD1Hn3InjWpFFXNl7ZXqUC/LatIn2NkxoUwXjXuj9/R
0x2UENdvNHYQ/jsqImb0O9QARAJl7zO5Q/z2eKLLQebwqEehz7ufedBGDSpmDdAn
6lX6vKPTkAoJkWi6t7Dkc1FmKBIvjRoX+LRG8di11IVMMnWdQFd572ahL8qWUfy3
PkooIFWZkulfyTaZCS6pP+rYkfzalTfJW3e0zH4yCbhUPoEJX9m6oNs3v1EUAJ88
I/DyuD9OlDfDE7kES+FjzRpFVCXrw5R4hS+HkUHqzGn1cb7PCXbm+fRiLdwHA0vq
JP1rVpDWhiCTILhtNqbZlT72Hr+t9ifDgy4zhvNtXwsvEe5msCdVQX3qDx+axtbp
OmYoqmZfDjJ5jB9WIlcN+U6P+QC6FH3aR6FeAKMTgyRNntwGzR7sOwoaOG1WHUp7
zN3LorMU89yFWUfXrvdu/QowMmale58WDUrY4n5VFYudA8B2oCQm06SJo99JRROX
9OiCFCUVRJZsIl5uF9GJnMRWL5JD8WgQ23M+lJEW5Sw/h9FOOEeWg/C+V/w8Rrj4
5YJxDDOdlAos1BYGe60u9Nh5czXEcJ/Bhz8wcYbm6FptTMLwspgq0nNhLaw8KOTe
kXeuJ+xN23dT2AMNnpdi/aguRGVXWF7+FfS1+SODkdar8qdsWlEG+jIrXHEVdcCt
OH8RrI7csS0abI9B4JOgoSS0IkYuqKziPztpdRRyL50ZDp0deKMGpO+pachIXljH
QmcA7VVu9CmbANAXh5Wkk96+W5RbipKnD8TjXFzdYvx1RdsI6JUVAlYK6IFLnSgn
ZWL9R7dMBh8GvmSJJg/lteX5pLkBtAM/6Ka9bNNTdRK9gUijEyubzjp/FTcM4rZt
f91o/kivuGVzVQPHBxGZJASlo8emP+TgVP/X3lIYSTL7euIRsMmypArJGrr3BmfC
WgR5hf1tV6HhGcc2KEsgGb1zSAg+RHP9damqrCF0Y4C20a2qrVScdy7Ymom1IObI
an19E0bFmOScoLounQomyWgn6E00RzS9QUHLzEIOb1ggWTQRUHzmBRfHZdZsQIdS
3CBGCdPK1+abGc5vXGe4bmeDynp11g4sragdqZaGmfmv/oLqbuUYKWBC3aHWZbyG
80cLrL1gCSCBtvFW2tWshJ7f61jHDf9/tK9m+rII5QxPdYqFc1TavJadz+GDQxiK
Ia3QtUkojY/0EH/H6Z03zSbItXflVhuThBZMJ3xbD2zcBr8KC73E8qC9IQuiWxKm
6A6BH10jEk6iYthnJuuCPn3cmxMzX7KOWS7jL1IDoWyIH0ofBeuIyjmtXSBpcLFJ
2kuE8C691kSkJ7Bg3BMZ17nw97qC3M+plg2V2e1930urTOHWtfvfbWBqttcCaQI1
i//eeiOCXBxEJOi3xYXkbkQDiefSg1ral027m2EESlC/sAJkffmAeDH+lIR3e+4H
Kaos1SdUcdsvn/7YrMkh57EYY1EO1Dy+kwZ3IyY+cqwXWvHdiY9Q/uYaGqDNT4iv
Hgw3MxhmufecXgaqRMpWcYgEuKqRob+nA3wrBSsRnvVQ01DWiObEP6m+7mjZsx/p
pbWf/Kvl0dm0m5DEekX0umV5FdGLXJMigfspwAyIqJWe/A0k1DlA30PzHbMcLd0l
jYURgDhZDctuKENPNbo7RpYaExlvwuiBwjVf1TDzdP6mGT2PgmrSvYZXA/TwUa7U
n8aWqu5yCc7Gci4cUegojawzx5QGKqdDq0TzMKIs2IrgTwiB+BH/CNBBh4TghsF+
Bt7gg6ycTGPKup6G4EYDCywAJ4Qckz9t0GEmqBA3F7byP4/gphIhHceXGKrvSOWT
SJRnKiZFcVDrRr/vSKRok2xmAZ/IV9TISdMLfRSLMwPwEObO58D4vBauT76rdmbk
pvKnbjckRFDp/qPlDwB2cHomM43ie01tpx5bIAVz/EWvMP03sxpRREE+NVJn1qR4
4NOSx/1E82x65EpI/P09mYjhO+4gVEwgDvL36kqR7i0va/Nixn1x7bowUlKCKc9t
AKy3frareZcsYjdBV7na3HtRB4WSO+fCrXZXZi2u8zenxPTuOmRfyblPFiJDRRQz
TM3XUx38x2WUuSAQS0AClCL19YcCp+KNc1x/RwtgHJqyne1TD4u+D27/tqc3yngO
/a//xOjdVfk+38kSxW+FlC3YTc0Jt3yjBRwW08HyDQKe72mcRQ4LSay97bTN9hRv
I0PhfuZmEsMENIIpNK6VeHwcHt7mq2GfuhvqsuWLoshVH1g9ZIyURuKayB/BwiNz
fCB/O17QZSwXLmRWuJ+/0YVOV2zbwDZ3KExiaV43Bgxugekf1HL2kbkBTViePfIk
E7ghweeRDCuWpSVCTw2qhyxtIFY+tEcbOQ9qzWyDKyE5lOKzqcedF1s1KrwIwAQG
DYs3FYfL7nbv5ECCs6WfhGd9hiKq5g7fX/7oaGQGzyasrDS+7kYeQHWhfZdInJMc
jEbKCAHSthUAYKf2Z8m2mSQ6ORFpKE71Q6qzjHsxbNBsed2EDtRFQrCqhQ5jUXgA
27iTTFu2YWctGAmjm3nlUQnRVSlDsmXY3JGYWSLWgaObROn/TAm36krSXpt4yylv
Uc0HDMOyo/2z0yVvmd/MXQD8AbRraMfm23Tp4jlplCuAZelTV7gJ1PDnHbR7acet
wPAUYzgakrt6YY+hxO+0p809yVhFAS+NFOOX9FoUCud7G5TkOwd7DDjE+A5ZrRch
e/oG2gGmp0j2bctd6oFwRYLOE/2RtKkmSjE92SXLg7kX4Tk5uj/srk+jULWwbVBg
c5ST96mDeLCR8PUQKRilHjVb6uq6lqm6z24ZrRgyr3iR5VqONhritoDFwn4BhLxw
w3OGV/jmJuj0O7aqJZNoBbwy0PgqUe8c1bSYpgCH+w/G28bmR0Z5FRkM/Gwm+eDo
+bn6hcthe4ux73tkr12Z4qsLuHst4DJVqMo27yfDY78PzlXPfZnl21M8DtiHd4Wu
lus46FgcLxlp5hIwvDRt8hv+oGclOM3b0qoVsVkrmv8pyVVfhxxWqWpovVX/d9kt
i2lev4e2xSGZ7s74TOj/knpqBIVQIf/64Py9cf6zHWKUlamE4jOOIXhxKOOIvo+G
PuDgaFULoifm0F7iSPvrA/CHooN5iH+dAVzOG9Q9e6Jxov8z1r19gQ2vGbBKFlw9
0PUKj7o3WhRN8uH1zzOoN54oC7Sx6zNRQ84bJO8mSTwKBU/LQZoc4u4Ks5Y3ZBfF
k++AN5UFwGRt/g336+0V5z5RV0PATJx7RZmg45TWYNgjlhUodCQasG4KQnsv3Wn/
EIpmiTjqX3Ne3FOv8NtVJc5GScv0gqUI8w7+vKmARchXFeNfg5fZiDavP1U6ovOa
J8veTXdnUh8+dY0hIDNcrDkFIZ6npNYk9zsAfgMssbhLa/Z2U/v1VN9zEuhyUMbh
tQ4sFO0SzFHR1O081MPVHn2RYYn3NWd/0eagGumIAYp1m7ZoVpiC5rCbE+/WescU
t5tv4vZdgYVVgK2jV4syxHsb8KF5r2QZTzhAD/CX12Ex7UFZLRKuyNPyXsZBVVyW
Ynjc8UKg9c1Ob9yFpT3GcYxIMd21jvs5xEmoC8lLYixoKYvKdXbnVwZ0FDXv8vWZ
WtH1uBNyNirAjoYsCZZxekrpf07P/ckn0xuuQDvJLZeSyQu7mvnR2FMBlrk21rVT
Ff4mrt8dwfgZ+NftTbEIRy2tuBXeb2Qah8zVxyP0g9+rhfbX7rLG5VAJiBER3oRo
yciEPJEHOtpg+sFwlwMgx/cjEmU+4C5EEx+OxYdRCa5s4sS8QqxT/vh1shad1JG5
HsGbIJ/jw5OuBIJIsSHl7uFa6fICYp49gE1ySEMEVysoimJhPtsCZ9RvEfsYLNoK
xxyAm57EWUocpg5BccyvFZpVIC2XmYIHkuQhDpqJgCpTGv0YmAywX7KAWyk5cuQ8
BUMQjiIn032RBK7iHAr7jlpOd6OqNJZrElGkXZJ3493xDatBv7dy67MyeGKNJQl8
pIVUdjWXHpk+ZGQVs5zq5n2oWtaMj+D8HbiegnKCAEUcR82fSdvodYw1+49ICnTj
TJLpixoPyv5uo3ozS7zM4/dn8IA5ZiNRwz2Nk4OKvVersgyZ7EtwJAHgM1Kc4W8W
jOVnmfEvlimZEnoqu+3UQWGMtbm/hmmSsq+xk5stNrW3kOo3olVWAc61Az24Md0H
ABXRrvlDDas9J8FB72AWfXv0Uw62nvjGHTEAqGbAw72KWArmQqUlktuGckxx1Ovc
ra7buFBlMxndFzm403wqORyB0n7HqvJ+4vpWBMew52ib0lxSH16K6t2huvh9pGls
W0kUWeVFWbkmYS0LUqzuoWlRzd4voGryIZX/b1PDDJONsKwL++PFI+R5peMqi1u9
SHY2SHDVq+7bnN7D73JmddJpdyyWtQ5Dh99H0lqB6J/jXGw9lvHcUlABkO41PdCg
JmqaNX0QCgCBs0HO4p3YsXsgFPOC2/x6GZGUQfcpn7SJtLq3IRPqWEF/QZwVWLuC
xnUKHMR7AT3W+3MY2d5RDI2rnr37EyOUoX1GHVPoCvDIORwfXOs+e308o/oZTihk
TJjOKlglMbbajGNB/p7Ktg+aliG1QtXc3wXmYX0uztvpR+rIMkKsETGrzH7kx8U0
AfZaXlW1w0WKjMT0UaQWulpDROGdJHEaYffHz5AYDQExmgTzVX0PY1ozudCYcIDH
xiZNUpDK0s8kUa47Dlp4w84q1ELutGkL70bikQrTNW+UvL2sSLWwZ9PxIrTn1yEC
v4uLCyG3T5pLkFOukw4oBgDY09dIBOXHMlqsHHQW+a3f4VHMCVQzZzAQKiy/N9j2
4/y3Wcc90Rquq5tWh1vqHQOaDprm+O6TWqdAtlLL2reUthrtcl3UBUWJUFNRsP0w
mM1J6c3gT86tcPnSP2soQw203hH0P9GE5HvWC+7kbzwXdtqNP8Yv/fK12+JXq/S3
N9IhKpNCJLYE7V6jkvt+NQBZRtq857ezlfoSxZGU2/lsjnK8ZtfIF/6Rrmeznr94
RZVJZH3nKUcZCx7yYvIjHhkDOiRRdFEHJt65MVhT4vK6TO7OP4d099vp6jyCpxRi
OXxY5zB+IR58GbX9cqjfW8Y436llBAQ7RE7IrUA3qW2L+In8Qubh2vzz9eLIXB/y
+cAV3gPb4oa0Axt5DG7yMeD3FsK1sYJslQFAY+Vo+koou1dQNb3I1hcd3F74tKbB
eDWuKXEEPnjU2GZnAA8341yFXFMLFhS/vkPynPUvGnlnHJz/N3EW+E/TNd7YQpXf
/gfQsTg4YVFtmY0HlnvqaWZjPaDRgPOeGrAUC+aYCo3AeVoMSMDBWW955aM1lAJ3
Awz2sYQOgiVMfXyxOI+v6yjCguNw3ZS+lYbsvb0lzlINgblhc+VDdGqT27YNNXcU
IxcUQNoEMfF5lyFH5CXqJIWjcgBu1dGwdiJt2P6GRWFHN8nnavvFId9ZySLODCM/
if+Yvn1SRIyK/yAK41EpgE+597KPoH++jXHV78qwICuygIVDiqXlvXpB2+3s/kdL
1LIlnjJzE4DBXK54BLC1n4v4N+vXdtJUnDD30rhXQ74dIuDbbLamwJ0G5InV7nQN
Pulfy5oShS59Egy1EUYgD8T/SGY6Klf4MXDhLYGCI0UwsvzQu7n5UZHU2ahDYkqi
f3BSyGmk0xhuFqIagWGuyOUFenXMMnm8UD9SsdMC4fijT/40SqXS+iExl/JjPjP7
+0+FKcP+U+W6B6a9BVAdQK1pcgmsWOPd7a3dmeuNNz4RVCNlkgHEygC4RYAowkKo
GeG10EbLKUNnjDM+zf113o3PUXYJLbH2Gbc4MwOqoCIsQTRmuSLIaueF6uum2BAM
4DGvsInLYEkhjIKSTSi2a1A7DvYmud7bHGp53PODH54siRhoSyPiyXK2tVEsZDzw
pRVfw43231srxkjpQMy208lAE0B18WRbTX0RIs4pAwJsnA9PvGOB0rNK9+byIFdI
vQ63i+cB2JPn0EScT5M6PFb8NiXmYhGH4BllbPTj+LRKrclFAyVWDCMJMrnQktpZ
S6YFI6zyucinQdQb/bJqNu0KhnHJxfqKpidKG/RhDAo52blAN50zEZCEsN2mMBPi
pjmIyOipHHCWsv3xz6Ih8rFO8yeJ8yjSdoDGSvwGgipG06J9L5c2IjCDoi4m0OOc
52bNxCeTuNvqfxc3tG6Q8yqJAsc2Q/XAzvGbiX+O875kpBXFjO7s+Bo01R5p2ODt
CUOMhX/H115uymTGAoM3Xh81YIu8hsfRpX/PIc7hZ6PF7gOcyDLix7iBZc+9pmE8
UrQHARWcnmIA1P7/AZxIrt1WWujyC3XncJC/eZGJ05cs83I/lCj+54PtdKH6ryCk
5N5eoRavmrn06QuI/1dd1Vf/O/v81dc1gACBCyxtXfHIA2/Nn4mbsPrmGi/JkhKT
l/QraKdl4ouDfpEZ3v86hFgJydfYp1d+dIPdlhQxQCun46MSFvFTnTJ0YApxk5Da
PYcbgko07I2kI2F5a5tKGFnFtI4NkYFhp7k3REAZALvcBgs3fzUUxb6UDGdPQ3zq
egJEvzIjndp7VwMOMBX9Prrn5TBNR2EuuBKbXZdjBoEvsJqFMkeReBOV/ymY8/zD
ZQCe2mM/J5F1vdfLiL/uYulH3XuT29FrhiIh9ebSvi/3l47kD76gzS7NzSIECuEl
9g1yL+UzNFFUFIlUNw9yd5xFGYQn95lchbCwHhZixEPur+VKHnJBLv++knASwbxu
dkur/NG5FIW5ydTWvcM99+ciigRR3F6NY3WWHqZogFQs2672jWhTXK5TdBRtGPMo
F3quVZF3P7II53HrQrqPWXwqaRP2PpKJln+fa2j6zhhfJArYdDggtXzmU9Z+TJQa
7RwAbYN34rZuqnYuaXldELMSp3dmxc/X9poUOoE2xJuBV5hFaeDqk64p94aB/IyS
F0Z5iOBpI0axKh/khj4fcHZ0ILxAa08uDUKv1Ze3E/iz0+iqUzomKAyu4562P9D4
PlhQhN3o9k0KjCmz8bgEcCvJrO7FxDqpphmDYYPYlHzGCDDlnrj30pNzl9opP3Cd
PVOxlp2rxCYRuHCe93wEPFGJX0ANrLSiNMX/tMbBtbts46ihlbpZ5hF4uJjmxe9u
CuSd2tNFOa+yuOX0rR9fdVi6Z39BwD7UyCcS6ZdPjPcTJ48i9ycVeMPyO/VpdXex
XgcB0EhhtJb1jAH6/GCHLh4Nl8L9ylRWd2utzoUvriJM09nI5UsOAqJz2cX4jou7
PVIRjSiA/HhywPn6HBelemVgzvxJ0QizalwadGYl9J3KUyM7QWhTjVWP25Oeq8d2
SugezdDOrBO8xllZ0ImEJygVqdJn/2BPvG/y9dWknypJgEpjfEYkcy6gmoXN+bH3
h8Yaa7xcoZCHajjs0nCo/JjHKtONDa7iZTnDlO0wDpn6zARjxNSjvrhd9YtVQLFN
kSKNOFqxthkQmpkx3Us0D/WH7DwgunGFNsodBH4A0e0q/timBIPh3hALO4dkPsY/
a17c2Lfob1pSGf8Ha2Zg4h0aQTwlODHsRNsHwsFVM4X6yN5J+THtrTQI8JxzWs35
haROFPfOP+6TOXmBcffy/mh/JJ89LUlG7oEyEFzJiPalFeBo2mWc9abblSIVQaok
5hEvTK1WVf3xccp+9B5eqEbPItJkScx1WfrS94XFoxwu5BoEwQUCJX76bgpUXB/h
HKqvI5n7VCrq3xPvafcFVpy0iN7ZylYNflArb7IwXBuWov2t8AGFN7G6unskyhm9
/YgMb52BtwQtM35KqmQIM7hw28wN5CEcv8PZuVYTrVQLE4HtSdfrO27hyAzp/Ojg
oGnbb6rju+Tfjp7bPhuF5693hhxU3jEAO0gv+BOLAXAQl/AAOC19U3qhomkv8EAw
nosQ/EU+WuEfuRlY8mdj2zTEdJwGT5pHMsPLTT5l3W/jsF7Q2BxZwQx1B+ihfOWr
1cjhQlZ0wHz4yn97GnjDGvVIG2lqJm1pcfsmWio0KENRfrVFJglK9KjUP1yQHDwR
qXbnCUSMqKi+i1Tb46PvENX8mSBXTQRwFjNj+1clY/x5AgmArz08eyerWsMqFkhM
7pc1JxfFJ9Imrmc1k9HEaJZKBh+nqxirxMaxdnRIg1oO3P8cG0C92HjCkK3BkwBR
ZyU0mPC4cAqfWQYKmLAfEOgLY0uiEEd1K3zq4N/x7uJdvhtJQI66BmP8+UTomfOf
D5DwdTT/cPTJmpF2jp4IhGaiajm3xZ/B4p29o3bYwtUSXfRy4pPPhY35G3X6eUa0
J/PqgqJmCGsW4PxGJDPXcldfDNskxZrjx+3PZNpSc0JtUn1Sv05CagkjsP+6TbjQ
TDb058fNAP9gONq/GmB9LUIBI+DcaJgdP7Om7hpAyeEzjBuCU0zO3Kx1Sdvi8/PD
VwMXZcPYdbVDcCrZUYxHMKf/KhBieDxByyMQplG0Ejr2nU5DjowOS41zWnq1ge/o
WthGZ4POyquwruuNNI9qi7XzRb2Rrl/T8xG3yezMu4jAvZ8V34p0+XuVCEG2LJnK
9tyLbMCQhR07TS/I8gv8HsVnBU1jhse14tao6iLkPD8ovIyLzL4lPWN/TX492ENz
LG90dt0beJ7rr7l54PoldznrCElILoGEht5DsR8OGK7DurGYu+/oGDYFyspFhcQ+
rujFUkXtmYcfI4KCdOfy5UK25AtIyjrdkOhja0zW7CQlSgXSNgNf28IFaXLUy18U
fUy04vNkDU0IbODJf/GzNtqJKm0StfvbyPc1Y+wjFxoWEZngVnFSH8VG/nWTQQ0+
vzMJdeTc3wyK6Z7eNt2m3Qvk3yXe7TklMMbYFi0YFlr4gCY/vZhlyhgmhl821Nb+
Cd5wm1+Ltk8Vtj9fjjJ/j8VMtztTrqg8r3qqtBu2RL94SCHxDa4Uvc7yB0EmRY/b
+SNnPYhOjM7+iOlpR8/azb79/O/24wBp/KrMBmH26ByOlX1HI1SzzIn1kjADqSp9
cGBaJHvKCff+5FT9xnnAmWJFMVmtaiT3Ogtk4oTAfHEDil6I3PSsbd9OzURSpgYE
A5D91VMhtOygQsC5Qovt5RQbCL00pxK33Ob79/6NanUllOBAe2Xn9SG4IM0UUepx
bRfRAeaBvhc9PjbnKxQYBSwi+dROCYy1cvLtzRy9lmyrDhljvPlxe0LXYlHsUFAF
I/VaTeab6q2i94gO0Po4JINhHjlmBPJ7hGZ21LLgudTO7QkkOxZ6XI761as1RqUM
owb0e6pC30PSuza73cClBZmDWHEzXqKX8+Mi1KtqqIfrWWqMMk9jKnwibuRLFuyQ
XebfYaUEr+5jHySaIG1e912iBNPXrwj39T7caV6nfLpca4lwHTb5XDAMD0OWIpho
d1ifqyG8qcEnLG8sCWmqbfprpQRAHdbxl1yo63hWoi4svmSkngvA8qQTjFacrvch
G95ig4uoAiHFuqkunTVmOdYktTFlFuedKpoMlffPZ8oZBWZBP17krB3wva6bGtBd
f+pmVK1vvaj3M7yd7TkmawYEjoAUlHlMdXNg6MJ8ODwkG3It8utp3k4bKAeJPrs2
RpD/s4YrpmFxvkmPieClkqdAdqV8hScVg8H0pPitxy3pfD31u+nDjcdzZuDEsZlt
xN36g2yrXnJ+7x8OBxJAzLAsY54ar+iIQ+3AGCAcbTajlAKZ4IApiuj7iLL6VK9H
dcaoKR6f+mBCqGfxt+FQ9sYsxSZ8EMzhRqNjiL3rDqT7iC/ZJg4x9C7V4JHpS5Ec
4EcvX80StCtgO365BACxAK79RUX+zpCt+JjcGQKoQXMVj5bXMJfJ9SnzHZOQx1Eo
F0LIjDIQPcieb6c+KzRxBaTX+VItJQIUAj9/ogkBNUrJRivZll5lbSXaAK8yT4aS
1M92WSC0AkkZ5lDAybeKbHIX436WuIAN0SF7W9Tq69KkUZkQPT7iAumgeE+t0Y6I
j0DBZk82xAC4OodSsG5UM2YmtNAGfNx3UCRnodnk9r9amWR4oTXuYopEUKSg4wp6
zj8in9PTf24Xcw2WnkuSIN5dAx+rILkY//53gpbv4hhOMLC5Rclkv+iR8NjdS7jP
swQjBrwnCdZvdZUyfm7iGe38Gqgg27A9L34zMQa39OeCpMbbBCQNKsaFQqQD4t4/
hGI5czcM0MP87I00Qz6DoNiHIhdXna2D5Rq8NEEZLoxbjB/O581n/FPJzzw8XcEQ
Ao5jY0i9r7eENhR/k6FLU6dqMEKKJa9ok10looz4vlisXq5T9rbSZ+C2enOY8kKS
M+RJNYgqMqbu7oo2oBoL41TPPIj2SU3drMjHEdLehcZ+clDzlkrBz9b3ML7RsvLW
r5jkuV/FFXza9OvDyfbPv5oIBOU5sKQQAA/GKcOUeRvqCbSkBkjS2/1xXcyEneS7
PORzpJnABIEl9j1aN7UNNXiw2ZSQFu+fiy2nqcFMS79Fh7ABq71wIMDZbNMyqMe9
013RRefkGj3RDIwZmFu0RHOxK4M9jCJPfzZ0PZ2oeXzVfi/TGQ//tVzboQDumxod
vG3s56pxDJB8iY9BcJe/qWzHHRwni8gB9AZDlJLOYnqeRyJAxSJaz3SHz/uo6900
aL/kOv8AANxpvXH8sXD3suj5oSjW9CaJ5Dw1UK6evAyQMIfks8Qs8zik0wnm6rHA
XFUewPXVITRM2a7XyflDRo5tQeuwEhXKqPlVpWbsmVlnFpl2wbGolB9lp8pBgnm4
KkfsEX/1zFbiVJLRUQkebPRB+98MM39jNnr0qIh7XOnFoAWj0t+O0WTLNH5GZxw3
TEow01ZtHp/DrsI4fDa1Hc3SYyR3jTNsNLfb2Hk9CAERV60VLbWeCom0U9Hk81MY
LQshRIEWjaHHANiQ9sB6YKTK8fl1+HGWyglXBMWZ+jRtw5G4e7pBl2Pk34t81BYP
PIYfZuiWuuTa8FTiz3dy/WMmGRJAabziRIgGsUpjRunpcaMyC/+9cNJeNjVmmR4T
vK2REdZ7U+ocpTQQzqkCjjW1mUxTpfZ+aaYmreO4BPgeIBdH7w8CpQ7G0ZqhOksy
E7cNsJyrOXHK8W90sMtrOZajh37pEKaTJEbxwoRTrsx2VAyRvt4ucaQNVdejCQgP
EvAsZHne4v35nQjDcJflAZJEHQ2Z056yinBf9Ai2okeYF34tYZH84OxKx3bLH+ST
+PgVrYGBOwpLwnhqsgeQOztZnCRiI89C/JEO7GQz0zqGLx7eSsIHmaQxHsR49VdX
ucS1lZRqWyIcgsUOG1M2dcAiniAI4pChfC/z2AwgDIRm6QZxuiCxEaXbHcLr+lV9
RHCbgSFTL2SmdywexqlEZBLgf4XoilKVXjioZVSNrEpJo6XtWfJTgJJmWvNYEgqT
U44Ma8U0S62ueTT1LTdWvz0zV2xAgFZ/DYFNhv2Davydj9HWc7ya/VJAIGHMWYUk
JuzqQ17WVYm2inZedS+Kk8C2p5maLbudgKepkVCyPZ9YyY7Uk0SQicysrv6oJEn9
0wzYKd/Y5FMBqugEi+z1IS7nye2dG1MceY96ZOpaf5ue6YXOzudd172gBzYgK00a
3XRDgHtNA4Z11jCfI5KjPuW98s6NzqY2UgIC1LFpJPTPa02YxcVTvlXdRBIMfACc
3LNUNi7dlvDtOep/0nypE92dc9qQwWvVjQmxAs5pGizipObia2C1rzRVWjHrwDjh
8J9bMQDGlEVEW06e2OAOe759ucNNECOTdzE1UrQw9nECIxmXHY5vZ1X/sDSzMXMI
7DX84Ba1Fta1LFtseDeqf69dJ/YhjrOhoOLyovdQK3VjY8dcx3+KFOkkeqiMHpV1
4KU7u1JVJIJw/CRlqeQLiwPmQL+JMMJDUFKvrLKpV2eyo6TXtefCBHb47+WPfcrv
IJQ+b2Zga2GywoxN4KIpMENT4GKxSxKEAVzmbsFynQ0r/Kc3cdkQeOD742dRihxh
G3XIJuB8c5g/1rxCeiBiulm/jBEV/ckanAPamHAYYXRxATGxWnpOuUISvAuMh2aX
mHs9GuMXG/Ihk4bodAk5GVj2hsrXtK/COXIXYqb8ysTszoSXmUqyBw8vn/j5K49L
X3Rol4ocZNiwOmpPGHDGlPN5aTv6CkudOR4QOaVBtaQNZZKwoF12+/xWEnCQAcgB
hCsLAEFfLAe28csyJGyOAif0mFBMACMUxbx/lVk8fKLD1GukDrOf9fXXQne7QYWt
8s0jE9SAo6gDeoPPfVbzsURRn8dPC4xuOrwg9fZXWRa/ZhBsTkrbvFaE0pfpl2X9
yVKv6RpIlnHAc3WM/TtCQt3HLWg84Bzn/U2esU9WoXEIyQtGYSBvNQju3ZfE8Na+
VWlVqqIY9pasQmWKQu/nLldpiBF3yNJK2vk5JK/y5sWh7p+JUo+nEJy9EjnESM7T
Ba2Iy+rT1DKAe78hdnDyMdKXfs8sP9RsYQCvbCexY1GqMli1LDXXCMwAq5FefMeH
FJ2gxC4PeC+agOUmBhBBK/qvRYeokO5ngwG2kuPz5lqbaVG+ivoQhtFxigQCjps1
6ags4S1oZmmyh+9USgdbb+jOS3koe8i6SWtqGgOOTJeSUZEPg6n2m6V6TnP3HQ10
AtZT4oC6iMJdvDFPN7y1DIl+bvZ+vuErydxt9wV7af+aG0xSTDVJncqflCExc/72
v9FGKPAiH0e2241tzqQJHRtxIw4UmsS5k9Rd2a1ORvMk7wYVVV/4UqQSGIElK5sB
4/hEVv7z9AEdrw4SkYFNyM3g43cSMAtQGbdY3gCaWeRaJhEy9z7yz3d7Fbd5eCmm
teF1SrFO6TnJFwpH+fCL5ScWGiteT1C0zhnZ2dVC/9tR132SzXKvHisjgq5WSxdE
jI7jc7rhvK3LUlK6RHyLhBZegUqh2WaqzhKQUNPjqsdjV4mBUxaY54GZF/PrS//p
pau/ZBJ0o3PAnC8ZC1dPRxxNzRTmyUUB6rwwxTUdJRF2++QgTp3hSPeWKK4UY71D
2q8Lu2V0mMM9+tfBuPmrJx4fmZRR6A0Kfk9gPgla9iV8Woh1DpTa688pTMrf7vsW
2tOW2+t/SDifDn8Nk1BzLhsVGlXdf5jwbwzK6JeW2WNI2hMsEo4Qom3DZAMdAQm2
2iV0X4IYbvLvFpq16K4lGGifONOGejoG163TRqHUmelYcs849f2reKnp9tAwE8dI
G0frSLwFHxG+DG1yEc02nVpbEKsk4i+wVGWznFrt3u1sgjKGFw+ONByDQ9zc4lc3
WIkLsa/Re+nVBr/87/Wuc/17rzDzD6ZW/id1nKQRwZ/HUdOfzDhQOkCxdqZddlrl
wd1UDCawk0+KTYlEqbxY2/10pP3xAet89MfSYMTahA2l7iMJ1uFQfW1H0mCYHkLi
NklQ1eXcdbn2RuBaQvkV+D4Mhu6lTzQNR2pSq0rWdY74mFLc6u/9+5aTGe/7OP50
E9p9davUkFMzMFs3ratI9vB6WihRgKdF2MpnCarBrqgi3h3a5u5C81PeMjkaYzxP
uqfY1peERfcDGmzCioYKRyyjNu+1/kNw6rM/RB2dU4s4S2B95T+3NZ0wuJC+WFRE
lrtWZvziIHIcP6L0YxI7SwjLLQU4aAdsur5GyZkJgTdNmjh0yj/sA2LvHoOzY8wf
84uLt/ZfPvrDva6PZxUm3mwiOczR0vD3t20nlYL3txfxhi8bpYFr62Af30RMUjTZ
7nfhtYQJ/9u0RCwf5BdT56eqH6OGI4TjMFhiE6YoYfsoXyHo8AIX0fSch5VCPp/C
rI7wSwseFqI3A8QtWl/8UX/+GvW+0N4k0l/4ekZ9+KsLrdmc8HRwEyygY5Nw3n9O
b+habKv7rB9TZt/0+iN36n78hvqPsxujw1VcPzXTck6cRY2LyWhuBwLZEvAmasdV
q4XIVnauGFLNGizwxTHtti/Iw0NAjUrNROpcV+emAScp9sWcCsEmBfKn0fRvFR27
KYzjwHjk2ZdpYR0TDr0cQCP+A58powc6zz4chFPnt9PgaANhKFtVkQ9XD+JfqDfH
G8P030C/Eft/9T9zCgJmxN1fevg8Fiqc58nScyoAoctQFDD8WyhZmU9KiW5R/yQU
37ECcQSzTowum2GkoQ8qU7hz8L8lV46QZfDSOJxn+RgF4OfyayzKsGJ+qA8RPB/K
lbqhsdP5NnfUu7PSEDqJnd8Fxzy+6dBAIchXJXRkv3kknYlxj5H5DVtu6YpuzXrD
xk9DtpsvfJGJ4o+/MoXsWy59QwVYDHzriakSXN6Bvq5/x0j2nqPPMSSZgmdCxAsS
PMjMZueEh7rE9FxqZ2Zzcqx1e47kMPwWKtVKurDTCWNTQOME2gfomiiJYvGNxJ4w
c5fWH/cCKEx6V9PNlOf6PcSk+5FsWXiydTBnLB/Y9BX8737KYCGtYGSjbNeFCB7a
ClHtwJ0LaXhngC8NWiEPMdo3afssPBup0LMIfer9JEOphEoC2AaURGB7DGp+3XKa
lKVlM2bX+IINAaQyNtvALeG/2kkQRdGRxyJRCtWQ+eXgdEBC5yPKW8T7sc9xSxHR
v42YGwOZLvM0Ym835KveiA4aw797hlFcbqxKEcuXxaH7p/m1Vd8gxyi9OWus1MKV
2Awop7YXVZT1Ta9xf8yy+QeQhFpG4jS4cPrK+DygKG1zhhSJ7aXFqMaeTcoO/uiH
AjHdnx5YMeyLEPXBEL2/dc6CGE9I1dhLT0yQFf9RCJo8aKHydSHYXx1MKUzlYukC
t9hDewBEVPKsyVR5toRNIL2L5NY6bBgDF4H+4ePPMm5XZsSnozL5987OhS5jncuT
GMN+9QTa3H/tcU9odyCIVNryeCp1am80Fc6/LYLUhmAlGDCl5nbAx1zXYuUvuRcO
trHq3QYCAv7KIT79rT5QCltYCWh/RXKVWnmTvUB6JgaVlu8RFK2OAEccDChF8Bky
+pYAuSF678sDrQ6sagsK4QkzeJ/7wN48ZGcu1AbMNcen5RAvWW6FioxgDtDPVj2x
VqTnuHRvwKkVy4MLESDQ/wpj9w/An3NlQTH2WvV1tCYu9/g2wmKSwl1OPmbsTqdQ
pkTpW48sYHGu/Qq63DuUYEhVS7vuxDwdNeYCCHi5UZNK+etP08Rnuf7dF9lnYFUQ
T+mNGYaH5PML+SBr3Ab0nDKLzt+goqeeppWAibUf52VbGuegvE5Ci2C0YdvVl2iw
b+xR8zLT9ayTfRZWLcyKWwMFbEvF2tty1762uI8FuTpFuL27x0VUjMOLNzVSWKFp
1nwgh7ygFIUSY2UN4yddITqb760r5gvpCIbKr6GYpUtrUdQ0We+DwxZKIek7zVlD
gFm1ahpP4ZT9b6oX+wWqX/AmQhOew8rImo1tiv5jlYJpDQ93d6pBYqsN7m9xLC8D
CxhpewtOQnQPNKNvG6S3IQP2HSjmOCDN5Z2UZYMbiQOFhpjRZmQzZy0MWO75PsC9
hHJqgLmZGM54zScW3Rs3KhUzDAZqTsbRDp9Vwd6fdaUnOCydikjk6s0kMZ7J07ja
UmxYytJvltWec/BLmEE55bq9AH7KLuXoAgdtOMjJRlYl0qnHYiqQVLLt7q1kMC+s
553NiMtj5GZyE1SKjP6MK7JYUCaf7+EmTmwAHmaC4wuQrrI1dMIxVcEkfd1u0eKY
8mknv+fqFCrB/+Gp8HVJcBHxgyu1maA3A2AlMuxhEgk/CUW7tUq3fRAYcEQqIdKx
m3jof72gbHuzOENeYgineXITXwJ7JQtleJXDFJ+o3+U3PV/2i/+/0xuOC14kh5U9
OPPxOW+DyOQAwRYZORYrDtZsY/cTqVAkYgxLvhXTxvNwLnQH7obi/wy+wZumniPJ
zf2wg9NdreVb+p7MImvOFZQzlSKZ0JetIfKOcqA/3zAs+gDqOy0asON+FB36dTEC
JuFRGbNj5U5dtxdTTK7ISk2XTrcUhlSd9AR0Kk12vvRYPJKij1iFrDX3Yz8Gdc1A
cE+J3tAEzMRzcry/FoVrHvbPSRqYD/TS0NdGdS4SJIMTKbdHxCUTrUJRak92o/E9
mvaJv6uzaLrxrnxrvRgunhk9rNP3aZgFe/cVKkoL7+C41xC4jhyn3gUCgyP3zA1K
D46gp7/pVfAHRbfG+o0iD5+ANt9/4brPy/KAA1V6xBi5qfBc2yQQjFy0+dCkSVFE
0zmBZddTUsYNWgDQow1AyrXDH7TH5b746up3deVMntpNYhj9XTkpFHFRzwbhRgep
n6mL7MQdAIM4YmVm7rm8HGkIHzgqXzGbVabC3sDvHw4omI9IElt+cYy0Jt0yiG+a
FpU4mRAZMvWvMG0hwk99h6R5Ovjavh6DK8kCcEwm4TZZ1oZzr8jgeDiPtKs/xcqK
7XF1Pu16dNlo37JZ0sQgLVCIbw8bO0BYIGr9/e+zkrhx1p/Igeo71XMkPyvFCI97
rncQFcbMe8D3RLUXR4lOA1eDdPURx74FjDWqvPfUZtHAQqbwraEySMmeigDV53ka
gAPEY7X3Mr7XJBVuu5jQWVi8iNW67gV+b0K+jh/7K194OeQ1m7qFv8sG1nzjovKX
j7SAteG/jDOvsH/S5F56Be9kenMkp8dmkoQ1vXT/hdgN5VDiIQqiHxqrDQoyhDzY
cnuypgMgb0z578PdkvDeaDPUcrET+/Mb1U3RE6mx1lQHRdk9OR1L066zORaiYSi2
BrAyHBoG8jbH2QdY/sET6Ialwkjib2I4hZ8pVK4DvfqSAA1mB2fQqjHQaPoBkd1Q
uNjsVF+ZP/45hjG6Ufi7YvKjWZW43qhRg7FPe58OxH5sEh7lI0xAyMAFszZGLJXq
hBouj+yRko/dVqSliw6HbJ3FpQWSYefqUy397XsjMnC6HcriP1LNz3m2VnRjfGvx
ofOV2X0Wh5zG1mipS+gHtZ2aUMTp/OXWTy7fHDYGs7qwWeyyv76ZZGnDZxF+80jp
JutTUG3fLRyPGYOV5nH3gNmhYnUmzvXehYJ7kqssowMIU5dyoJdfwMBooNr2psd1
TAOgEpddyg5Ojq9Y0bR2pAHL5EvwFz7yMC2ZSVhyrZ69aAUaRCHzKQ/RS+T5vtmJ
q33ZZamrtFtVuGYu3+K9fgd6W/Otb6tZJ5kY93MXe2qASjf6pFNfEE1vyPLVfgG+
9oKCX+O/p91+dvGD/zIyEmjofWCFyl8HwQSiJDCSrMjYYaYd1hbcM3evjrOz9EmE
nk0YCIRg/XUT2MKsab8YAGNZtkJgXHsQCyfFBwGy4GymEbP5KDi7/BjFsZCk4T2v
KgKjuWVwHIkphXSiZqh+qdT6bi2Y+iC6lmYzHVjg+cvaCqnsji7YvVmCT6fDuvXF
Hd6QYjxGBIJJbJ4aam267g6T96yawVqB0fh88/UNtcpWpzDTXfdtfMU0VNHujFeF
V21op5OdPmGK/jYey4MCs0j9aMK0cAXKP94yQwMdUg1EvFhqfFzDQMVCIYwe+VI/
gfeV05f4dFZz0i8UXY9ZlzATVGJTvgd0knDfXiDlsQvGtEJBwKGC8mpNWO3SXVAI
8z2bpsIbdc0GM3id06ufAKw9XBVXmXmCsUe8LURNgq8upLMSfvS2RXTLFTVLCj7l
ss4QQOG+tVS2MNHx+/0AxAiNivqIP6ZD29mDJzoLVojuLDTy3a1VuqDvF583Qhjg
dXUwqywbMS4IUOfU2fXaojC3lxmREOPqwvd0vk2+vQNq8m+LPPhKunyQuwgpE5i8
Sqquzt285POGmLPJzJ6ZnebMCO6+STkG9ZluETjUOy/XbzHt8imaLalDs2T4+0vO
cDRyMiN0WY2J79ByFBmy0jk/75tAZbQFPa9PcYOK9pHbJ2m5hZYp6LpJf5nRxgnx
Y+wHhCMFk5Lh6nwDMuBAVe76SP+IeQ3PuZ/JIH5ZGkQWXdYkEutbEw9NJ2QKmqAz
tv3aPhmalB9nliD5YGoNLGrfKPKQwEIbSfKlsZxcY3esB8xFQNACTtHkO3UcjtlZ
BaBJYp57gyM6zoaSXg3/xegUUYO8cihHVgzOT69pmKuruklABcQkdBKmX8pOLtPH
S2UHKi24kbMsowrOqoQ4/6tAwRI+3ZCFeGnaiZEoDTl2TMwfzV8fRh5RJbcJ8TOx
dIP9m10Z/YtdzMtWRlC8dKdoUQCuoNeFRoDiHKkWMX/gZZtzqNEJFlRDt0aameo7
u0e0lb8sKDyOzipTNkQbIX4bcLyXbp4Sw65SXAL2tDUjHDACE0EyTT5LfWSiUgrZ
oN1rGZUh0wvr37cqGM2YKBhk+T4SxiPGNbJ2luNn190LGXw0Pb6mUEy7piVIRRjJ
+S8TKYLD0zE6B2jIcjwK2yPeLxQQ/Hg2dYkYR34aAhPZmg5CqRHvrZ0UvTxC3/in
gKFw3zaeidHKBHvBsNGj95ysGRFox7S3OFiJzb3IIzrSuvVmLaqyaDV4rPurqi69
ziPJZCTJrvwHtFBtlZ295vJ8+9Ons5LCr2ArT5paDPLSLQJi9JzLZZJBJXhO6sHk
gQNbaqQoSdRsQS9g/08+znoDZDsLfqE+it/5V0bFUn4eoLIBsaRKKrbKCHPoLTvf
bgOzX0ljnAM7ZGBvYtvPY8CgowNjYzfz0Fq0X15kya8EsaP8hzey6yVi14U0Ggv1
TM7Rnpch9rUy2XDF9K9+qVcJ00dLDLlp8q+J7KPCjfptr4iBImxU/PaoAKFA0KZb
cVtIP3ZIk4VNHqI2WD1YoIBqn43SUMdZrxDCgnYs/T1+q7dAKMt+6d6OKVz8naDj
ewyus8sgRveMWV9WO7yygBzdJteJ1zSGx5RCQotxHvfQkmxjpQoK2kscwN5jFyJl
9ewboUZWKGE3kZLNG3BQKK6NxqMAr4Np1Yx+EcqEgK/JIbq7x5lj+lPhLgMGOICk
Qr3eQkdXy+px5KJxmGmR6/JMvsxm54Fl+IJA8L/C64JS1PwgO90NX7K9CgNVfSnL
D/xpCvoJyNK7wNwJipJM3v961zkgPHAZahKd+2+1iCOQLu0eKc2FnK2EU6l1uyqF
wryfnZ6mTG0Pytl8h6RebbgxHTajc2pUi18CoRJC+M52MF6+h7FWUXxCHjuCQMje
ETCelxo/+Rsdbsvb4abmRNwdffpPLj4S49SVs9MNYnWKc3lWYkAX8SAHEuoNJR10
5mKJdPk9SAh2hzKD0VAVNmQw5zqHsho93fvxymbAgoLcvb2MlUp5nvUV+eJdYwjj
I8GyEptXSgLdH0rXo2v3/zVhqlhHossqyBKF4rDPWKLWaa3WqxFduzOgoInXUA6W
znzb5XmCYrCL51m8gpbWmQL38GpueRt5WPE4ar9ajLr30TR0ATIPOww/f5UQsX44
gw4KaBAuRIbrXk43aqLtfUXEv5skEOA7GFhN54BPp5kx694BCIkZvLuHHF26hWG8
krqVBs/mMJrBz6MJIPne2EuEci9J4KCWl4biT+HuzLECLViK5dEEYJxsYu/vPdaY
aeuXAPRQ/25O/eW9TArTyfDVGcGD/mrqkAAVHgozsteqeYXy8uewPLm2RA3mm0xm
/Jg8DvlhWnriOFDuFhUJiZgjidYsVR7HljjgdvaCsWVMhXvljLS49lJrgEwVwu/Z
mpw1IWDvygNa1Dfj/uRbQR4duyymNCTl+BVJtUsQ5hU8FActtNVQb+lZYLIj5rrE
tyR1JDh01MXoXlXQCHVfUZq2so6vwXZ3KAQ5b2H8loKWs37QpB+qBY22GVKYZHL4
prBYc3OESOb1dmXEA+ONKpI+qPRMq7xVi2LnYKutEFR4stU+rPeQdrJGhMMn1Wnt
7q496AufTqVkJMjpiRRsJikqyZ5iTV9ktVnIk2vzUEgj98akLj8ZNKxiPRZIi/aj
Cx0cxaz4LMMw3rlhInIj8N3W4IZ87HPsLPZAe4aYJ3JlWmTFMZQaNzaUdnWFQySo
AzOUEwWQ1VdUpoWNPtDkn1B78Pu0BujoTBoCeZPIuhB6Du9Vk1406dudcKeYTP3Q
osEALoaMaUUgPQGN+re3ZBec5qapc+uhvL098MHvIQll2s2JvEckPBlmGB9+SKa0
EOMAs1KoCFB9fm6iknLP5/nPXwIIOrX1yZ2V+r/T4K5coyvUaesj+YYOtifIMEp7
SjQTwYgzPWaeTt15usnYYtOfcXkL7AJdLXBQ3THHOZJnTQ6blWxAYkbPx2J9QG45
e8ryNJBcIMoBBIlkFVXAOeNh+bfV0cznHNqWypjzjozCNMg3jySB0LNJdrhmhA/P
HdZ6uAC9++PdK2tIaKHwZf0VzIpbOfSFpVrxZ9kjnw6v/qpR8aPRUPVwfqpq2Rym
wTpUB+0DiiE/fQfkHgFmkVYBuEJP5AR1Oe5y07Q0lgqMrZd1yiJcGpt/gI2HWL5w
j8p58eFjkBzwpjhIsP46r1GZXgX9OnjH7pwqFcDunhgJMf1FJGsu/r6ouSSwiVG9
y7DnfNvvi8XPAeMkvzRvU1Zcdgh3PdFLrxXgb8lC7so57mke4W15OOVSiniNgN31
e3s8alvOb0MQ3512Fn7FkiunAlwsRxak8Oq5lp094bz/AN/Tg5CkYkCuWS+WNQph
68IRpg2ODNyzci3qHvHNvQbFzm2dTQH6UddJrLB9KXW5rZhL5tcEEa/ow90d9SeI
1gcOccel7Hcp972VBjkbS/RRxDPwD94QsW0StDW+6IBlRs8MnHpsQ+9grbNFoWl8
KmhSXTFU3u5zQ7YxPctFLREjTvApvBR7V3sk6pswwTiD0NsAG/pTFWWtGvFY7L7r
oiLxtZcGYiI39VrEZAHU6VDWE4cxsDrDaMor3mqoqGOaU5+aBbS/ZUzUXx2OuFSy
cuLV15yldMEjUjfnAQJynpYili2rj+GCr8N+feCtraSxOY156UjITlNXJOz0dBJl
YZJgFmVMklbTb6VVQgx3B7TH06rdRhbz4XNHX35qwra3yldlLw445fESd6tqYbB1
+QL/F3xFE9iHiMIF4oOV2nJxNB/iSAcRM9NT+UcNmYnz2iSFxWZilAzG19t9PQCu
5zhdynwRVfhYW09hmPFkOq/TI5/bGq1UjDP/ioFGbYoKFDBFtLjrhXVnZ7jXjfmq
38XSm39i12gEk+PuGfv0t15gEVz9AYA/ddeldMPKu3/lTWdp4tnr9drf9YDsc7AQ
QkWZMolATTrz9+4mFhMr1hEcjdfqc9PqBe5DPro3/KocY4UGL6H4pljFleuPiXvd
GuCWaGFDfwzjkwm0Ajz91Rv7D60Y2A6WBg4Wiflk8pfMoTP09UFDLtymkk5gbVDX
rycVo0wM9rdbBOsfYgteiH2++eejaCRJ5WZQASZfXQaEs3lJKhXS8MQa4OYYDAW3
xg/OqzNTLxQrFAiU1Z5DSLq1iEjhEg4bAL4rWlagveEqYg4+MgZtROa4IecEZjjK
hjC1fKxmZf+vUd8+9Cb8KB5oKagt+SKYICim5TqeUEQNzZsXrHPQpf1phBWOZH2k
M6e5fm8xnSNz+SDmtBuYjIZGDv2sE6UMsY+dYay4aA3N5AcTWYNXp8DQy/AkiogM
SEvVqV4JVOO+V2LWaFIes3QETAA6OO06aq/BTVofMv89Vj/StfdfqcdVxX2Jow7D
kPc/unk3WQGfWkLQyMaSXMtVlekRb2rQo6Dk0T3C1sKsLqo/q4Xh1VwjnGibkaSk
03sFplZ9N3U93u+I8PoVhhxcPRw4D1bbUKAUBOxcZVsqcenfVOklTi9+R4yuJFYE
MRCobu8zaEAoKpb/yc9j7tlEg0DnSr84Ax/y7P4jgEGh5ZzZ1tk3TcvfPdMvkl0X
lHWHzkTTgYZGUKxC4c8nq/C+JOY8bwfnw7jFPI1nFjncLjS6DEnfFgUq+eZ4byYY
4ecUiFMeLxkvnOwcPNluwJd5MJmlDkkhu2mRBW0aosorwn1fgGecKDATHhVPWQDz
hCZdBh7Es+XMyVlC9DGfjcN5sMhkphkKttiu4PdwR5RwyXxXPb7srUdot8e4CabO
KZNfQ+tvQ0PyP8x0k2tfuPOEyrx5rKF+5A8AH/+j+6QNfZNBSC2pnzX0PpOK+iKs
ACRqaAb8yo5d9EPyr/qTxuSVMZd8S0h13KeLBXA8aypJOV3jWV3l1fM3LEVL8w3a
FBRm3U0TSYgfoGbgg5MThBwao2UmcuhuYSmVfCY8QJnhBJsJ5JN8FlHLelt1w2SO
5YhLDulI/7LvufUoznRjFfB7cK3FbSz3sayRngTcG9mA5ZWwOBYBF5yFbvJ90nSy
8HA4PbCAyevGlTZBPqEY6SEz1qTX5clLXjR1qxa4GcvOpoAIFz4iYQuAGYlNUo9o
K1V38uqEhMqsm8+eFES+zdNhaO3oK37ge1MkPgykZ0PhWgi2ynrN/M2uUX9ZBKOk
mYP1bGwr7om01kYNDnehjimuE8Nt14eLOGyMRhNY69EZ9JH6RCpHrRTGd075KoDk
BubdhMjOnJJpxTEtDU7kN1X66yvjvw060C/UecmhGXwqj3qYjJDgARh1MgiDgPKL
Dg3hHu8FRNI6DzfZ6wzCGBpVGhn2UOcXp+jNkuSB8+8sM+fmHDNDfKlRQLy814JO
hS5qhRsWkHwPuInmG4EW++8BksajIn0Sh8zxsNRpZUeeSTx5VPVEv2weMGZ2QJLk
6QLiKBsgYaEtBS4hvozSietb+Urtu8NeU4y9k9EFt7DeOLByjc7Io5w/K5AXunLy
EoeFQ7llN0Sexal85g3OfIXTnbgtwKfOiygvusr5y4yrp91KUR6j00rrRmViZ5k3
6OfSBmA4McDRXC8UPXorNh2xY7uRCRU3yMNd32uhPwEMr/RpHN+e9a7xKkgxDXCn
T7JYSTl/ykmChTrCh6h3ujd/PB4OPeZhu5CO77Y0LfhO0gMGxqimjLvfuM5v5OET
LF0JOhSOoPU5Hj0ZGRaVQhFdRPjuvuS5M9t8Uas8NaFuefPvUZtDxbxcVWtwwiIt
Km4j09nm6oqL4cRPQvzXVcWXjV8XoPNbqY+DZuyvr7TDh6AIxjjsHUOT6Q4kk5Gu
liS264k1VynErKLNRh/l81g/WHXmCdQi43wQAdC9h/tgIHDLcJv8JKsAFXkeSLIL
5Sv3EHwvCvJuYQFu27NUHdMsC0wt5FtyHxKjQ/nGrUgHbzYIyhsrFeNJOKW6yZA+
6018XfKrY4KCk3lWeye3ThWnvbd526JoHIDxUtAArvDADU7m2BsBYfdfEW6jWPbP
0fSXLqsz5DbW88XXba9XRcrR81kStpRjMMb5cjZzkF6okxBriwN2bkDrh2khyfNe
h3XK/DgZTeYKZh2ABsR4INrvybwnbdfjK0ey4BQxJKWyl+XUUCvypGIl2+r4b80h
Nq3Bicvuzp0PAiGTLL+ZpowgXRu0DRh8HGrRiMhAgB+1uUYsImtE9OhYiifTZ7Fk
LCU4eiTuSq/dXfZHkfNhZN5yF3RK97yV6nYfmA90wWhIR8Ikoj0XJvYyvvAAVYix
qKi49UuucKtkCU0jjBOeSmHKRUFWVu1wS2hdU9YS3No+0d+d7OxFonro2CYL4981
XEsQb5Xj9joErXKygZyM6ohmrqoFWCLlxAoiW0Vp39FjEGWq3f8nmkIfu8QzArlz
S/fqW+jdQmglWYms7GZp0+VGAavleaAQs71v94f0ywTgpe1SYrI/RJ50oRmhdotn
fz4XYiNglCr24SBhFAJOQsQmp83KIUBFkFLaGVIEOaEqsFFxyZzi6pyL1et4YynA
tNuj+gD0gXM93DItNpkJtIvnBWhwbB4VlN4RxlfmwlIgLPSPLqJzcxZcmKAO/pLj
uEYAieyH9hvLtqMkyjHpRz9/3Gtb+12lZJNKxA05lCtVQ8HjJ+TzcJ8T+onL5zAg
Ecf738mDteteC6rZvAgAIFBrOecuWxgT+HVNIE+IsTX6+KAA7HtHH+N5G+DqaxCP
8vzDFtxqH9lOAfNeDqUwA7WUiYSrWesSG30IHSvQGeKJM+5hAgczDrVRYsSkFTc+
u2DAupUJ6amLw6gcnFphb4piLyReiuzQWmxJ32jUoPoK+vSh4sigvC5OXI7DK1QI
Q8JdeSD+LsjBL/kEW4JvtFRv6xtWCMKzTWKT8DljBAoLP876u39yBxzQeup8Digb
ZpqEbjotqMCQFQOJMkDLLztUPT/aYqaMf/XiGc54x9BsJVmYXKS/7J6fN1A/4nXB
gte7g+Uo+YEgw7R5gtnGcy3YOO+uNmvOkuv3VqpZ6Du5rJl7QXc7Fb2gtzzz7Bnb
X7TbYtNDU3SlELYuKu2yfLijV5QFG96Ns3J9MtbYMlehv4tgqFxR7t+jOP2FGt6O
SDfI1M6wiq2lAQZZcanv8YGF1oe5LCMeQShjCFAR6OOCWrXFGYb01HeMJerZdORz
NihQoz1sq22bzdLIPpJZZJaY0pZtLmS6iCvnvEF0e6l2FlsMaOuOZ7nyVxzXklKr
mJ4NRLdOCBw9EvkJ8u3m/mBl8/o0jNAfIK6JyG6/8r9B35ANuFx5BqkCZmq1KvCP
dodW5cAuhf3qJmrZmh/8UPLLd+67lW/SwJZjCdSo6W0Is/GbjKqeZJwJR2BVUZQt
VoJy6AZrUnd7t97nO62CA11c+b8/SV8nlDq+kdUV7oj73170bSlMhHYKdc5YctTX
zo+9hjuD7JXl7HidgVoLRfM8CVIyXyJJEN81dt/zPcEpcwPLEe621QGhcbJI2EbG
Wzzpz/zFAqAOxOa2AjYAe5Q+q5d9tufXzn4GzUS+M5HO48trcPHaqDqw5g2HPIB9
/N/Ot544F0IYFoalSZLypQclbf0kGLGJgMs+wv72MfOABW0KNzYuEdkb/5SCUQtG
prfNHeh2/DQ0WaEhpq3zYLMxXnguiMTMpiUILBLj/4lEzR63g78Rc68Bs/KfpNNb
+8aB3od7sOXqYTS9dQA9uEF+DRhY6ogHzEecUCUAlP75+JXcD4UCLfSxZEQ1JJAW
hcJe7vrBukG3mEhcdicc7J1vmfhIDdHXNJmauxigqSAuG9rKsAOxRNGunD7r6F5m
jW1SuZztPON6UCBoSbvt2IFe2sh2RJ17RE+X3lrLU97U2CqFKmfiNXSuHZvrwmYo
7OfkD8Ximd2xg+m1oegx660T+pUXBlPCL4/X8JCMKezCLCLe0J4JAErvg09Zxeax
Ws5oC6F9cW0/mNP9apcyrdiZdi+SZpOtijXL8Yy3lpfHIarPK3DFNL+5zbRKO8FI
7pgHjDkbRw1s/T7cdkg20lUKXalSwmO/TXqHSZYCq4mICbVjQ1nmnYwjL+4rek+Y
SXgREn7ZVrC1yz0r9FWH43XjXHXIweGoX9sdNftKHj+GKezEci5GgybPKGHbGxmR
vYZk7dQEOYkWnz47xjea3pZI8Rhx/RshrG3YMyBhd3C532oJBWl0wxNpTdBj3Wxi
iLSvo8n7DyAnso0aw+WppFR/4kiuU0Cs4GmyqJz6BXhIBryp0qHxtuRn6KC5UDIf
TgvxIdWVZOqctaQvxsC4p+7XcaOXSvcRj8vaKUU2J/7lnXYEVnXVHLsKnIjgFloD
oTpBrcsSPyZjwovownw9rUFTC9l1g0DSyKbs24rnXbPWNocRCd/j8ZVXPFeY4lvv
AT8q8OwhXW4ctSaVsXiRI6hHbMvQqQUwdr7/FDz8gl7vnn6NMj9HX0kHQT/PN8yj
nK14ydSQYmIbrQtYINFvlaAfOhOBAmIAf62x5RNtCcTDeXDeSlUiJSA4GQgWa1AK
eUEckRPRhRxV8292H96CJmFlFHOYj1jHHbKJV3N+nDUux3LFbd22wrfT/QZzpw8w
YXBVA+5eTXg7AfPiHpF3MMjewaKWawx86GzjH19f+/FEaN8lVlmGtbptRq4x+pL2
sM4v6MrF3JKFReTt4xABSf+JmlkqEtvFi9E48K4onYTXtcRc6ILg1KRAKGTBgqIY
L11t2oSVvKMmBlfkdfKXxsqS+vl5i9Pw/1a1/c/GkX2Vx+jQcYyz/5ZyXF+2lVmG
VaFWwy+oVIUg2HmHjTWIRn3yQjTwGuSugnA2vlpuzQI2LXf7k5Vun0TEArJVo8vp
yQzO3L/g9Cvmzd2nzHb7vz3fktA10zAbHOI11cnl7WG35+dYvVYpPPXDZfhltzIy
EogNUQNWDhZKDebAs0HKifoazW2Olcq4rKDgkAxgMPAWDXQCgOhocx+p5zWdSjHp
QWvHUAtli1zHeZVbWclV1oSbClzd4jkU7qmIN7Wpdm6xqXKpkrwyKaSOj2iSha5h
LGdqySSRIaymATvCA5n0Uf8dKHoCrqMeoYJEbBY7yIRzprOwsgt22WR9FfAam9LL
LhHh9p5xgN0EUao19vvXSo4Am/N6WXrcQo1K9l+EdKghUYnrAMp0PoPWX3jSu2wk
Pm3qbMD28LPl9OUZiRj/eL5Sw/deped65MDxtCAp5pwxt1DLeC60Ceg0KImXHJDL
K4Yyr6DpaIJwESuOTu+SuMmHcIjoYwr1ia2wfxEbPLsWZpEf5mWv0/A7oEfpJXiG
wNerwwWaVZP0bA9mszUyJHdpl8zxg+QC2zpu7zRfVB/J57gDN2iC7GmR4YOEjhrc
/pKO8JabPK2F8As9yVdAYzl42316Dvw0e+x+gEeMvrBidrnHpr9HYdWRhKNo4mZU
ifywvljp4R0UeuyAtAx5KWGVDBT72V8cCKPTSHkBBd2lZd4b8Qe8Eml+HCcnr3r9
yJhaSrOdxqZ3fe/nhn6gh5UHife1CZ0fLng2uZdj3nL3AZdNV4VNPjO1QUnS9RRG
l9zA5E/phTtk5GNUHdtswPFZE6lxvpQIoB8phW74m4Hz6n5Ny1OplE7AZxekjdRG
O9lHjU+MuHA7M4Lnhg/hT3FVqrQXJuohkkzvZ4/r9Os839yBohp3bIFp30/GcUbW
kRb3G71EIfev9fDIXc0BCGlgSUjrrdguPMzx6OhSPOQoYuAauZBSxZPJWOU+Gcs5
puw4omRSdKwHQ0T7sVYDx92NrGZNuXKBprnK8hTWfnQfyzyrtaf3hDIolL7M89C8
xc0YlQcsVb7UoGiEwG+8DOHZR5nCgtgSoFDC8yaawUPYJjWA0ejkHBozXv4PxduO
dYeOSwvT4EQW2AC8cE+C2YrjElw+PPeh+XYShRkuyU/kuv+5l8SBvRF9U6wiKzUu
6V5AchTVoQsVbSrQQAJKvxDYuwkW12zdaouHe6wH/+x8gBPyDYwj2fWPY+8BC/L2
55NMcX9ph6pe++AhPLoSN0vhl3CYt1lFGgc0CtoMvx65oA4f3b6wJhEa9bGT5AyD
LqtCnuAKekbYTZONShexZUCzK4TQJBi9mJ1qpm9Ayv8P/86kzkZa1Jm8vz7KufGt
Xqw/6Z6fMDzSMQz9xdY0XLD3qzCZa2IYE44elmQPOXiYnkBnDxcQQC4GioyDyebf
Fu9EytrypXOcDDp52vWgGLPfhmVSVGxvemCaDOGeH2gZRklIcmZLwtjidliAXE5g
RVjGRWBIMkJnvNFD/nD8HG84k1o+Zhtb5FdnA7xUaECP1YKsTMfCWm20bghi8cJP
Bw05sJum/X2wN5KSrTVZWFG4XaNGUyu0330ohmh8+W+Cie0RUrsJtBkdeeGifW3K
+MQ3yxuiL4sKLSD7E9BpCL37MuI6EvlcDxDvYB9J/pzMVrx03tnXKRNYYKvW+Zm4
Yo1htiwJD19KdBRvmcTixSlWqZ4JzFKBl0WtJEqu7NGH0ENKkURCNES4Ol51kejc
yUVYGYkq4N+0KI+TfC1ZVEwDB7efh7frFIHxb6jSFHIi8GBIuQOtipJOvHdKZwan
f+ipAyQrwNKD02oO+kn5SB0J3icPhGLgTxcwvM5R1EAJLDUGaSkty3SRoGn+W7x9
PyK6CpWsPuE0nzYMQha2QZeTugmWTfpcy1HGKgbyib1/U/O804RnB/AOSZax3lTX
vzhjKEZUmHGkqw0cAOyuwSEbX7D8NIBQtlRSr3URNvvrgRcexb3f4HkgLt2yoHVh
+fPPAYWuRPZN6mOz12WzZ7Pf7k8fP0vv/sUvkoPKytd9u+cy5qDZHuIJ2dAtdzRZ
x7+AoLyHKzkAN60LwZ77uQ009yq29EVd7yiXOhdM5vlIvQwW+9mNfD/I7AEp8pks
Pdbl1YUVfS0n22tIQ56IjkVUGGbK/k10pk3UN0OZtkPKX7c/nc0j/EYuMho+Wbst
yRI9yrHT0xfK0ouYP+U82GFzUpODTeVgqvzExMmsy1oDfuj/+zG7QZ16Y2V1VOAn
Ri30V/8iGY1bMyxFDKfdyS0PqiG8ey5RNJABeaLsAGpGLDr7RLmUU8dOAbfaP8Vh
r/RwF1nZdJ7kiJtBBLcNZtB+9MhaUhNolt0bAOqgnmh62Uqut2mnfFSnXuVIL1RI
+wEGrtDxDroqn2oQLvfVBjJl/FlFaQMbuG3dE4qV+VxCBsaZ8Z17Aisv7OCEucFs
TEmQJyArZikcPljIstt2Z/IxE2bdWWZdLTdxZ+GSMJFwdi7t07AuYXyxhKGjVK8p
j+HuYQleslfHKVTxp8AqAhZwbauLhko8NazUH6TuW+34MH1l45Gf7wsfX9+o3Idj
LeM26bnZ+GPgzRf1Qld190p+fFYwSkCV8wNrtuih/fOjy4RnRGJC0R2vFb24yAvN
xt0J/5QOowe6gz8lMAsCAVXg7pb8QiPay7AebLe7nPUKVLt5GRZTvWeap1qi3dFV
c0TiCnq3jUg31Ocqju0hhVw1nJKbvEWa4V/XuUL6EI1GWAUH2/NsqAx/uY99EKGS
PGb91ULwH1Z0baQQ4nb39xX31uXfCKMrZiikabBQlZirQKBsu6mxY2XWQ4paBIS+
EzaIY3kcdB6RfFyGh3H/nTCKq0z2Tb9oHw0HE1tBggofK2OWItR71+LWYUwGUDzc
lr2iH0o2HbN0U1Oaaxcf45l6a8p8u15TSbojm/3EmeCxS/NSxJVWQMR+bu7YNbrT
YztqgUxQ6O8RV07/bHOeeoQ33b7EFlbrgl3h2v/OBw8tXmXdaKN29MvYxxojx+bm
ZaIwX6DuGCTqq0qgNmGTaIVgilnXuE3TfDowvQhYe/c3toYlM9r0goUM6yub+WFc
1hmIZ0sYE//fNXgaIaDsoPgop7DjFJvQa/yDnCqQyLhKtXp9PBuaQpH6u/uu0mX6
M6mwo0nhYqM+/TAwUOWcjd9L8fIWetaNeRjdLOlNMC49uYTG+YE5AjbWRh6m94IJ
wk1YbTnRXFax71cR0azDrMbR1zAEChBukIMqQhaD8sZxRE5k5bDTuUh8TAdRjp15
qvQIAgUfrcbPYFgh0MfWOR3W90NkufjuQsKlpJilB9tyvxTN25S6VAM0MzbVQLpW
Rc3Mn5SWatb4LIO7CAwfHjsmdqhWO0Zy8Y25QCDrCq+b/3yFoeYm+FtkGD23s6jz
AUHj3k+27GbBJpQFCy8KubkfiQy7P8qywf9ygCDxWqNviMR1XFEuHlxOzhSqgTZj
QYIBNzbiSo3szw9D78g19cq1PVZYSfHXpeJkU56WyeFY2L1Q2FbbZskBcWAmuvGd
vZUozM7cyUQcru2pN7xGQVKkmRDxjMqGUF/Z0KLTZzs0nh7ipiQRfUy31+s4bXyy
KSPWR1Nzy0CuKHsrV678G6MpkDikjkyn5mD1SzYymk7oJK5vFz6bJ9P/8cXRgV9b
CzmoiedTn8S3Hzq9MGLieYh/8UailQPQjiDqrjZg++MoXMBYW94vZmL6OAXwMHyG
utLzXWvHm38slQMtAQ09coVOWYlUrA9x5WL1FPqichI7aX4e7YpqM/0TGU3KGv6q
y9XwMX1WjCNZTF8DQJ6T/FaEfB/oaWX4kPkX625lZzrGCgkTh7AnVT6wmqGJerPN
CWafB0owNVmGbJfab91bFDGlSdYDAXKzstAQmJW7PvCQ198wdOWeTZaCNbk8/nLq
y5VmKilKi4To5QolV/9HoN61Ti25fCzxfrq5wqI2QCe2mY4QcYy/GCkhJR5CCQtY
s8jrGUWtnELgPk8FPpzEV7GnSxRL7CP17DoJZ2sLJ+iU7yt13fPwunPWtenJ9HYs
H4Yve1N2BH7nnWu3VNeuy8zIVatbvjzbRIPlWKapyDajRJWPDIVLpyFuupBFVt5P
IFuOLRpDOdPvySmvBOsb0JHr5YWqx5GX9MugZCgunaDLg2cedBJRmGVB5DI6g3Cg
JZ0J2qjw4+VA3KC43cIzyATmaJI7q2WZJjR2dC1qq8bOvmnV269C1JUx5o0QAHdU
HMgGlcv1EmcMG69JO8RqUrqxVyGIZWQivT9CBlp8SLvlIWre3DSp8G4ZSCwyuIum
caE0ay2QOE7x81EPwqvQ98xiXz3Q+w3N5facxPDSGpklyb8Ko5A1y7bfA9X6DC5K
QfN/5xxE180eVoDbPURyU2gARsZR7i+NGJV4iHRwr1WpOQKTWsNFd+KhPo4Kx4eC
i8il1XJc/mXu8Bl2CvUr9jEu5ypWmuv+9Ng0P0HuxXBkXvmSRYh8JKwJ+CyFpuoP
0PxLTcCP/0l49EPtI8PF9wVEOuJCzVd7meJk8c4uyvUT1Ql9riM04ZVzbtP9//kQ
Wk5WZ0oNWWd7pd0LOzFRku0yt7HVKckfEQYDyyb+hNoRMqhv/pKsqz+xRV+VSfbE
AxGuKGbnygSE6sgU6X3cdr3s7wLDbDe0UFb2Frfl8CO7r+4pP9EtPdfoftd7ZeTw
HenCV+/Bler8tdSTsnsUQ2GX2H4v+K8W3XwbdcEh0ZimST+J8rlKaRGM+Qk5ld5L
UmFqUExQZh30JkZWDWMq2uYUkYPflKFeW9+IqesFowMGEHT+BnMkHi9n5HcHZpWx
6QGg7qCwfEVSIGrUGveAYhUZEa7DqBscYeSwE/mBdfmQRKegnmIDudK1c6ALGDGU
EicAanhlxgBNql2fikcY4mGcoQrEsL7crSRgdGltEczCDqxDEqFw3OjqNXzvrsLq
5zwthEtT8sBZst2tV5ggVzPOws8vbSrvlxCH64Th9Cw5PQ5HDfr4fBsVqToFwE1p
P9RI/RQSLFxQN3AIfLggbgSNnyrwP8LivNXuHsjGg4/cGqc4CdMXeOcGmMPKBAgM
gvhHbGGbTXC8TGjKm4S4QBqSkuUgJjL5FkIOuIq/VlwcSWXw3Uohu3uKYi0CKYXG
f/DD9IbjX1ykJZXjGZX1YnKZrsFN3qtI99w5KEWtBbkF3OAzzJ0ex+UcjotYSf4w
yLrVh5L27lSpB2AfaeR3pmHt3BUBvZQW2JtUoscpFyVy2gHvaRMElGfeHifRNhYY
Iw6EeYZLcctX7ZVUesGh9BHQ6ZUk4dujUSpMiQWu3qFZkw+iS8LUo7ZgV3zXlT8l
bkueBePL/USxfsjJ3C8sNquhdm23FtG/SwNhoOzomHuMZAOTAzgW2grH3f4jK5as
N3oERWLcKSTFPcCZ+e/Hgk9hoTK9lpTp4lQqlCzfsgQgG183yzpFkZo3h9uc0ak4
hJrtO1OTjN7bl72Mo1kyQAv8KjNCRVo7BQeaVS7qWc1hLl+j1lbPuPPeusXIqZ58
+Dgb/smTl/z04Gsl99PeaYgGDJD70Ts6xZ04JRHpkJiysuDWKKKHNRh/Wv8T53KA
x6vNFsIl5/rnytRIiWK0Vg7grtyk0+8gHJRCJvyaUy/4uBA4ML474tMDXBEeZeAm
vPSC/tNQaabbrUgfHrES1TGPjKfgbJtW/W+RZ5XdOi0lQt7tAgiKZ4MB5AFvYPiZ
+1KlSm5Y5osL5EUEhfy1hAxATfgnUgcuS/52+Y+ZswsMSbK1IlSBlckxnJlP7YGz
dyGytR7EYielwJjTPz/aMV+xfs7ZzXyMXqo0R5+1t90QBqUdAz1hSxpuTkP2/vPd
ulZeD78E6ai9dyPEBBASVpUwU38i76TSbeLcoN5fgcRon6tNjAvgdCpR3KVfiMON
ouZP44I9F8ql2hhCT+Xca0Ohl+/M1Iyri9va52oTTjPQmVIRP2Pm9hTe8+o33OvA
4mE+35Mbl0tuqremtAkhOdgPnst5OR/ZH4iuZPP1w0wnGM+rCQ/1GBFFNSodC7jl
dEUiaK7Ab09iAiGzgdyaf2R4ZUEPcSwbnPSMOO7hgwh22L6cE2ZPgcLlTOKNgwhR
kjvEOIM6ZQ3ko9XdPDZhhQ4gc6/R+/sGA21wkis9xM5nZakxqoVXzpj8XVn15RF3
Bfq1kfT33O5VThJHuWKuWQMQ+71XRtFf+7WXTh2QzhOQPVsc2Z7isfii+QEWk5/O
Rka4+yAlgWPL1Hz89tUP6kupAIe/byJni0clgX1OmPoEpuM8o+S1rHeXhZBPqZ8e
JBgkfLNw6LKUdyotTXo/Buzk0HkxRZaS+/OEWgfHa243pYm9Ez9ybC1qK1j4dOTq
7jucuo2mxbV0kQF/6JOAL1Y64UwFOgNBfrAQWZsjfKO3OAkSy7rZ9N4Z/mm7Khe8
9KzDSCJcYMqJI7zKSPsoaawsPQh2/lWYruWyURChOL/UnoWvaXhya2z55svPbTDS
OyhHdMOq/RysTpbkem8ooEpjnu9uz9gHr2U0A5HJRz7r0jQUAOoKkWGfzkmz/3Xx
MiQN3Lo6Efw2IeEGvogV99NrESl7++yivo74gjgKKMEnPPEaLgkJTvGbE1YRUepo
p1/4IBRNikXMOux/qd5+QjlRSX6Kc8ExVJwxF9QJYiPBP3Yhj16jxuZ19w4H8dsY
P93eYThwQ0/vhEFh3aC8e5sEFwcrxWtDae3HTKu0j8a0KJV4UEpwb9r+NjE7A0cg
AogqmSwwrQMNpGNdNaaGpIpKzqoURssTQR2oV9B9VobtEDzEUCviGhakHeC/mSl1
gBYvjcmElD/QWDQ+lrfojClMg7mdK22gPCJ5EYCy5FKyWX7W7Vn/iXkUKLNK9RN1
R3ij3t2qvaAQqrwSLOodTzQNmisOXVT9t4bJaLZnZQt4dTZTe5QCNyCl3gUbzWTS
ziPGpXdIr9VbRfL9lUm+85bcq4h3qtgoi2qK8SmYACVH9lq3L9cj1yxMtbYS4K1D
r8qFnBG1g1U9YM9AOG+pQvSl/0hWtxoF1fduM1N3bIMKYXnP0kRCrONBhaKgW317
82FbFPPlCVZ9t7v5XV3XeqAGruOwUbsuTaRzfcacmzR84mJ9YnbFm2OkyfLAcvj1
buBc3tMMcacYvxvRYJixQkbIcHEE9/IduKwvHciDbManIHGaE0Alw+pwO71pN945
e+E90CUA5IRdMdoI1Eyvl1yQoInII4S6NqXiruNPOQ4ecf4tX0VYnvU+jZw/0JxB
Ou2IXmd7vu09PNsyc3ogpWOO12QT91S+OKZaN44DXh6OZ8sMmaQoPblSxy3ShFnw
EmYIOqOQYlC8I433Xr3quRiHWlNPIOKJaf2WT+woJrQnJcK0/I4hA3Y5JkMbqyv/
b/eG6sfom+9/61lBWf8v5CY9Tc/hObZ6uUXQciQsmBbEiz7fUHCxQuWUwefte+Nz
2o841LRz6ETi5dNLblsCE79Nb4M3O8NoUApwOlv+j5/Vss2EwjJfOvWqqcNKYEBu
gNtzlQ+BBHqSUnRTXm4wfVU5MCz8ubtL7/ThY1YZfJ/R+F4Qs1zXgx9k3FmvWZ7E
zt9fkUY+pNQQWWYut3/Flcn4mXFn7pufKVDscJThbk086DSbbUtLhvpbbx/7fwP7
Un149WHkEBlug1xia7RCy6L457yWBUB6w9beYighNVJ2O9x1o/9dcAv5/ZKj1Qp3
z6sCfwOW8YLxWtuPvub/wRNXVDWon/vhj7XU2t6uQrnyC+hjPnDblU22Md8u7c1h
DJ+FHGhjr6efuqQl6BlWZ/wNvpbLOh2pvhbYk/Q87hBcizD/CZENpa0SIPomIzrg
o+ViV5reAS7LryeIa1N6uMve4PMAxrgIAURMvWxVMEDD0BhJ+Sa/5Q4HIenQf68l
4i4MxMSH2C6nOE6vP/CWdab5RkZNjPQc+G3leGSoN8jobbbKYji4O5UIFHle78kf
l8N10xMFsD8bnZZ/qg6ov3FJ0BS5ZO9K6HeUugljbWkNVgW4hg6z/YRVtgeUCApd
FKdXWDfYq8uizudBuqvkdPFG2mEuQbQVCgsozq516u9+szC9t+rFO8deruIUM6tM
9i1V4qpTa4PRhrwWh3omV0IyJdO5ZUeGd9EH3Nsxu/gYHK1AubkC/vJ2KtT8nlzs
bBls8BMSfKRkGrp45Jo5HDN+iho5x8Bg0ZTkUO92Q5bRl8Pu6YbElH4epx80wuFN
mCRMBzlTQYX/e4ot/5VaemDcWPYM62wj3ISCEfXCqglBmkIAEU1hzAB72W4FW7DS
qNbDY/sRVwhGkE+0UFSNTApxtfF0P2m5wLJ1USEiKtxAPGD0o8zRUM/LPYTKizPI
WXksj7uSUQOyCvvzsa24Nn5WBwqiZ30XPAFWpZZLQCasKX/K1Wx1Q3UIFEg2MmA0
1L/WWZ0KC/9FHKNBZ9lYIC4UfuZ5kBZZl4IKhorS4RV+nF/O2MeYgGMPDgAjXnVo
E0bnODojpsKESsysqyAYtjMfwkQVpMLrZMVH284atyQfJvjKUGTV1SYbmvOYNu+X
90iEHJX6aMRRF83ZdJVafMSgP29d9ARjEfYRRtTWfkeWYZc4J/9eRplzOdJVh3QV
XtMwygtMQngfy2ffG6ctDAvXc5YEknzr281OqvuefIpJtzUqdBXXagezJCiVKELd
WG2W/pyHcNkLKN142aA4v2/7wOw019MymVBReURbcvIvL8ocUJR7LG1qkgRUtB7Q
IjTNZWemhrnHWqXu8ZNcDqU09dCuKxk97ASYuMssD18D350v8/qK9REwDEu6qTMO
ic6FDJXjDvenfmTW1D3rtSL0BK1btsuvOsSTFHeBE5WuArNRwFxJYHc4GwA9Kugs
N4GkS3Pyr2hWsJwLTY8mwspUCaKr6CmE6x3Cd7hA0vDFO/jAJ6VvA6p+uBEsHzO3
OvfL9An5E6I+99W9zmeK/onTjgaXRWcDYn4eMZG7AdOGfY3mo/MqGJTUObWCw4F6
H3+pKShoZ3Ei2pMwpctbK0heI9c1y0DTZ1eWKmWqBvuBYv7puJYlxhA2apgn9aZS
RWTIHJrJLOAao8dBT14FjTV0ioNysjKcSLW2QeQaDftg+wwNirntYg93dY2ZMsfy
y4UNaXTfqJzaFb7QYIIVMIMgv1tuVSfItT5QLjhC0rrn+D/CT6YwSGxdAhlSMB4f
qCmeq3O5uzAz3GI/nKSUu02SYSbS4JHIGOwRMEcvi+haovpqWpfqRXSu56DAYNBl
GDeBcxPago96T8f91hlQ1xIL0gKC+mWhor5QRpAF5GXDUQt9g4Woe1RC3nxFbYni
7Q/A2PvuwDTagooGtijdTNA7+koEhM5KC66hMnlBUXq9GN94WMtwhiguXHIJAReL
YqFnZ5HEu5i7SWUH5f8hgH0NU2T2GfMrsyCeQwSojhbjP4/vhWLEwI05KWiQGAEm
z3uzE7ToqWhKfVUQ2rfs45SYt+HirC8F3k/XnUKZivTa3BCrI+jpxeOT48YxGWO+
Qf8+ITTUbzi/jN/qAlawnKehQr0DQeSQ5mqvmKDCK8W29YPmIamoU4HToLkF3jnn
g9+U66tX9/KvPnKR5a53ddfpL6pvHdKz25jlk8zpHnLSMR0BCKmpXj3deTLC+s6B
l8M/Gb1+VTF5kiRwyUhdZNcxrFoiRvk0VTMrfWbxfgLKQz+IfLhWV0Om6djxp7rh
acKIGUigUvubFlIiuWedg+1AdNePJPye9kWxSUnQhIdr2MmBS1vJJUH1R5BiljlP
O+O47HWpbSuQDmoZMbvpqoU9ev1d5SMJhtJygpBna6ieiij3jUJOO7dnj736QI8+
5vRJQkY3szujoOzPpMmvxBun7aVnl/J2Fae8TXWZ84dzDGi89lB10v+7JTxMXL8L
NmDWtlGSK2+rN9T1wE9PNLAg8Gfu5byu1CgyNoRHzfa5CioBrbNWdbfOO4qeJJQf
RxqlTpk+cBws74JBFdQc9fZc4Dm15hLZC7+97AcAX/L5lwu85rFDXWD0Es1hZka5
zNYYxYeo/U/NTuUPKuKRuTqmW179Gn1GZ/N5NPEa6B7Qx0fIWHWGR3O8OZY5GdYY
RubcgxfPBF2DkRC2pKJ/1oDQcjHQzLQYAXSLtsukYv0+QWYZOpXSv3WrgJ4LWc3E
rWyy0J7+O8FCRmaCDBONFLuy4obCy9u6bhnr9GaHQZidErBq62HEcRB2c9HP1ETV
GKXAmkEhZThejgsXuZLQdhpmvXIFxOBBPun+RaZbF6zrcC50G1WxOWe8jT2uBNEN
5ICmdsSB5jBatWhOqphR8wVZkMO3e+rEO1kEeBoQO4iVogXGg5fFJYDLygW/pr/i
oFrixuGJBcz+AUXfPUDD1RAoivud7/eCzbCX1hbY0eHAPcEBuqmVaB8WoXKLpIYv
Aym5/bqGjM/uzLS8Wr7OeKI76XEzzUirq5D7WtH0z1rhADsAC76AfNOLWefjVble
kyiRr3dln0Z26wZU4tkJwRgRmS0XiM4uzKLwdvWz/FeuVNVLKvJFrf/mCrT4N9l6
hmwpWJ7FPuPzuywOlopD/qxQoHZVPdxXo9O0Bw/gAXf/kbYFUZ93X2dDxyA1a4Jd
I7sPSe3ivGk+WWXPTW/aPHRSRdgYHHyQpis2Urjnd5fOeaBS9eVIdL3t7//FpB3P
oPoSq02G6HLYaF1bHTalMR5URRNZ4ZETNeEdRKmb4wg+n9/DJrl3t4gI4VZ7vIUQ
hkAhWGAR8wtORRPx03iv9g2mISy6FR0qxpg2DzTxsp63VfGNkhDcv3AvljxgxojM
iQC9ef2TFwAWuH2Ds7CEOz4K969VRsAw6iApHrQTQBToWTmddn2OcsUFVwpPP13Y
wbE8ZYYmRUpa1GcjhffPkHrQJWiB4u4qFo72L3wgkQzf87Hr4p8KBZxA2M2gxgBT
XVOEYsGXZiUUceFpAZ5nML6Be+bz4hYlZc71w0loeubVDv/9EX8A2vwVj+kp/PVD
IL3rUGg260PBtlrsaXuy7YpyCQdp7R3xnXMbe9bpdEfWyvKILUDY8iHDr+EnbqfY
f13b/BP8Ks67rcRAznwXWG3X8UjQ5MfhASi2CuMeZrFinsJ9tmZ/Qz0avLvL/dsA
xIfC/hL5OJ6KgdEbePNYJKPGgde/J5uH3zX0t34b+Q/APPIVZ5hgl2c2Uh6soa7x
Md+DKGbHs5WBTq5TNCgGk5sjPOI23V/oRsvz8W0hc+ePjLKfKCbkBdcSoF/eAXTY
fpNgDL41AMQX3MU4H9tdyAC53AOVaKG5lgFGIBsgkmN1b0Af4go/uAGWB7B88zrE
mnUDqpRni6XqmN8mZPkCs44FNCk6/H3fY3erMX8k/qzzGVFYY2yRna3rlGem1UVC
YfVLFdpsppNTDMrZpIodkwzxQ1tQf/2ozcRflj6Hz34+lhU2sbxavYNlRRQyb7qu
lqDmH5NmdhD/W4+R65rteJK3Ta1C3MbZOCe/nGkuKkgB+pB89/SnRs7OcaiNDzLj
IDdiG+qMkIJN03UVCK3+gdpWCY0TB5Xs9u+yqMZy7meKFGRpJ6lqIgFjlrvlDHl3
yf8Zku8yb97i5R44e7PeJVlTMcH2w/g0xLUDC/SP2IsRzZEsl5rISvIQDHZwK6SC
dnnDE3IR+sSMPHPV1JpITeoAovkdxGH4i+50mdUerxVq2YFCdp1txxEj1KLpbQyU
Rj5kqlvoEay68aOF+nOTPjS2bYJLWs+pFE/ArcMbAN2yHfy2HgnJbCeXoS6YndJY
qfBhh1VJozywWL5Y/1g3xw2zsgih65OPhibG6c0woZ+DZDJa1nSM/17n3bUPyudV
uQmLuqGQLN6919lohkn0X8n1E3/o1n54deNnUZcV6ERDDpcMVNldpwrvRq+CszRn
PU+GXLMdCIwo/2H1oo4XpTL/m2XUo9fC4CIsLuLnJTT3Zs6vzIMH3Yd0g9YI1kGC
7Oz4CnfJyWTS0OW+8Nqi+Ztei+sRU4QwkEqC1/HQ5W3Dj7zPylPjshlN4I2YxZOp
SeLS516xDojobS5IuX3/KApfytX1DIi3M+FTvsdjtaKOnUCDWUXgTUZMyM0+W+Ic
HYMLa3wOEwjSP/c2v3BYcgIINsSNS0AGmkD8KestP12p3lX6x8h8LIpvYW0gY+15
3KLTI06IKN3wQaJTPyh7XYt7c6ANnzZvepfz7GAbtWm+k40G0Y3rrGa3l1L7l9eM
4BEoonIGu3P5w0EB84Y7ubRdxRTTxltNn8n1vwJ0/FLj8ZUuDd+ANdvNjIu4puj5
AhlckOM7KJt0Zt2P6ry4TZn8co7ben0AvdtCQiaWmPrE5rN8d1syT8rtnPRRoz6S
YFBLCkM7BanTCANTVgYzUTPkeS/jdtIrb7dUF+bAWrovf/YE+UIl3QFouV5s8Zp5
2JutWnULsAgCy/WzcNjlE7Yd0pEm+6BMYDBJ4u0Fako6WI++pimTi6OBYH713a5T
j+sCXqb9CAdSwnBPRIebRh+AL3XTbuSmlsGmhaQLcGBygdqOpCeDXPfsTg7OVD67
i2ElHSQ/RTLxxCC14AyFAHwj/Gf88iQrOSpY5B1sGjk7mWcrUNF4q6be+Acj3aI2
GAkNm+xDt5T/7TPm8x1hLpw4X6FOCkaK5aJYKqAQeEMJXlNkWlIxa2a4s6naP70Z
sR1/BQuCw5cOPTdCGdPXs45ZAjWrAr0+Nk9jKwkqbdZ4NCmo6enxiAoSJ7aMnS1A
6zKPFkUtgEG0mryYu67EaOGptP8QgBVfzLdKsvwu0l/d9xitUZsCx66YHrsfZY2S
9T9ljRUh1E6duNbGaSqiOjgvsjR/t+CwoBWZAl5XupvPNE6krQ06mgVCpSJQZpvK
QCHSuv39/0Y3lxmVo2YwFKs+6Hcygbh8l+fTprx3UQ/X3wfQ2vJyoJD0gpqrbirD
OtYANiL4dS/J9Yw4cawjhlj5ZNb3KS3yJvGXOPKj1Oqp9GErZVqFn3NHeP/3N4X9
QrYlCyzE7O+Z816vA58uFaGJvWjOvf60ayRc202wk4RZNzMFHWNUMtMD7MfltTZl
MPnj5MYAfskrjqJzSUfmZpkN8NHVSdvSISHr5jqVOSw7Fh+tc/vTNOeJLxuOFgSB
Zi4flGIArN+0Tzl16nR5VX7yqaR9bB+xI9lb2l6CJ9hmR+2dBzASJZqVMsgkYr3p
lrwC5yRwvHuR/YwPhNXIYUIgyGw01ESLSptVZCaNPJLvD+QUF8CVXGFt2S2IiwHt
8cxqL8fvcbYmInCsyvnOXaf05hpiQmWXlmulzYwQqZKmC5w1XqhuunON6KhExJoV
rC7QP8Fmh6a1q/mt6fbAxCPqHkL+2t5OU6sa7buspO8yssQ4phQfvG5PnUKe2067
0L9dXEM/wABy4PYNIapeC407o7EyEBB58/p7x5DSBb1pqr/xL99b+tFuNEfUpbRp
IOugsMr0SXefUVXMLUslxnhbneMBBoaBQQkunrARXyIUqbkC2+vhZPUsZ75Nhq2V
wzqEvN+unWIqzpaTacskmFTHcuiBx4yi4mXt9sruBaa+5t6nNLeF9Pod4NLJvHur
dwgJ1uAZl3i0ZMZUU+56hHuLXojlf6J6D3FwugizOMIB+4ZDSnwupwBlQbOCuZ47
hWksv6E2uh8PnP6EERjbd2/CTGMspXN+eB2TASwX2+5JBTbYs5gIH9+NijpfID3t
y+1QjsyxofErNmU+oiELJLIjNP/1QN6Gr/YojvDeogYFWYSVfxaTPro0Yy6W/SlN
4ySyOKIhE2j8MJBLXNhRt/a9O235QnAqSKZLcKFdlF5nr/0YoeoulE7Pywc+4G9W
dZ52bxS0MS1CHCyMKznD23meGEB0U+kxLa4NCkCUDb1PUtKwrozj4DwwlX2K0hvh
oAh1D7rSx1sdU4+/QSfLKFPIl5s9Aj7+qpZQb7qGVGXqNUrwwInw/83uHbFIEy2f
m6lw05EOd6deFtv1YQzFIhI/QIH/kgJNtBqYEvS4FXiinC19t6CBPwwb+gWwSZIM
q52co0/WV7t96YS/McwoS5S0m1DT9i2kg4edlBmgBispl95fUSNxgKUUxZUydxw9
+ZLcC8DCmcoMzZoBNWKQ4tq2Te+kksiwlFtRQHdYbhyqMNLLVtQbItU6drIWWxat
lOS0S+WSZCZKR9/VmBVmD4vtb3IY7RxKiMxBa8zvycPAPnN3nUeoUgx7fpUkAbJo
l4ZoqpqDCGFb/lfM6C9RW3IoyoPRMBvOTj7Buwo2EwSQZYt2OTLaeWB7ALIu/l8O
N8KELkZPOlbGho0OZWO28JtBgHm59Ax/qRKmLJ7dU34I/70ExtvQgSIwFN2JioPM
cFe5W4D6OXPHi3cpc9lumtt2yc3VRk0Zej3St0OWFC0Vwiup7HdQ9fAxJqQp/vcr
uAXoIWMhYTzau0eyA1ui7FHpkECTPbR7Ve//2fj0AjX62fd4qu2pHbEf4BvyM3z6
/4qmC8vG/wl0B8PRWvbR8at1ZLkmVCo89rx3+SjpC/1SKDfyM0twSKIVaIVBvThP
mf5epHU/ELIa/DN/QR7reUj8fPoKPA7wbjsXpPZCmCm/c47EoHsn3x/2MlPvttOF
k+dWaS+XodpI4yeNXW7nJCGQ5go7lWUSbRF4Ddx3H9UJm783Brtoo5TrmNHoE8q1
Lpi9kNXBwA0S6ODWnvQTzE9OWgy1q8Jm1kb58+bht4Qf+C/AUxEe+rSVHiD6t6pt
/NP5lAyuB1ZlRrbRqjjzJqoY6nXM6Elb0ZwHBiBrMpDONmU0/wLh1s2J+CI+rY4u
ygQR6kOaS4YEPWc/vNIA7nRVmQnn38b9+lc2xv6dH9ZbRwuElYZ2vo81x45/E4BX
0Ako6QrC4lpGozIIUjjSu+lQGMDhFpo44jadcxNNGOqva4cQLs1xGdCMcma/1343
4r8XI/cwXD5kkdnbe+skU0S7vXZTWgYJMlrinv8V2h8BskH0tFaTzC03N6IQdkbk
Yag/J5mbsReGPG62XMIEncBKrM4W5xgTQ/CU+DU4e2BaLUKys6mqSLG1lRQNl3ZH
TdqxapnCwzuiwHBqZpzqhJk5fZzxnCm/J+sEFaFBGA1sw/98LKPMfmYDy0IHzy/R
bYBLY9az0z6CinBm1GFipYezFdkEon0KjArwnqnBbWGEzSIklBOS+BNx6d+0pGjn
vTVT5uFLASIaPqQtTza3rqMMB9n4wef+PzanBNRXrOG8/jCJTG2/n50nH9+MOeyu
gdpS7PeGxjvPMObYjz2VTleU6Mk5ULF9x3TX1bH1Vk8NtrrNeJpvzswOzLj6C67W
ZQDsvzoxjVq7oQdW4+CnF8QQidxDWenMeAHQl8qmBXGC++BTm4dOOIv0/KB9CaNz
yaXySqJT8wes4mRLZmL0jfG/7/wGFyPHwhBxIWXXw8PVhgY86PIsuvCbZCQKdgD/
imhSsTrgJsa0Lz2quKYeHjUGeEAZWeTxBInrZ/e0EDe9Gimtu6XaMS4N2ewYSS8T
BOAhTt7ueQA0Ph6WnepREVjq4aYycuwzYmZaVmDrpaB+mSEi9Ec5CvGHcuulAmOX
y+zhG2v/2rpKuYD/q6SAqDHSEJrCzoyurBcwKPyR1TiCy8sJI1LKYzZEc3Jc5HN6
080avS2TbEwDI7H9Ay1UcDkDJMqXKeY043kkKEjn5+p3KkEWHzkjdysteox2caEk
z2aaDb7wtfawDXPp4ZBD2PnHOy6M9jlVaRbGN/L1yqqewX3dWCE6FGZ6yCuuapDk
Jie34RePB402YjJOflRNFVXyDsBZV1/VZsWEsJWfUvTw60fYMNvdqppoYTMG66v+
QXTIf81OTwzJBiukfzbpUzVDnvV+y7QDoJp7eNmBgS7g2raYbhCy4+nRxZ7++y4w
q+2n/4wePCu17D2KrMeYxIbQ5LUqQnGlIPnJGNsVYz0eUCjgLDy8yv5suMsgQFOP
zKWdac5oW3e+PFI8IKURrr9i51D+IO3i/GE0ip8oNkD2uJlciwC/tfdK3p1HsnyE
4QoBKxdgnzWC4i48GbwgHPKhO1Rl+skeTV/91XCuka+eBjuiwdevACUW2MmC3VJF
FU3AkBpI4ZaUb+96E/XqkW9GCNofaWWOR0JhqfuhjbENF6FZOy7sDlN8/N+koKi9
RAQFNuUa9FSC7h2NZQfe92TVmAAY+NatSuOlsu4EwSJllHGG5TQDJbVJk2I5yjXz
z/UXHMslTui/QkJYI3rfYM9aFRjcZjgl0OGWifKM1xWIRPCyTiaA7usYxJZWwCka
PrN+cABRnjFHKx/f03ARIRRLFLHe5B3EzV/KyemZgOHCb4gkTdzHlJWOEnEO6sHl
quBzxpJaVmnbHISyYQMU68BXcSvPEE8aWqvBn7sA6g3TtjTsx14x+zZBlzBiNkTN
NauwrOv5F2FVJtutSs6YpalfkRJtxZd+O+yr9UZc89gVOo2ajSdnYwmqU39+GSkw
RfiJIwxfwNTR4jeXu6wU5CphVdRS2lWlwY3qdoX8h1FUm6kRdguE8QgHUs/oYhru
rBuebfd8AajlxFjJHSIPDh/jy54yMjNJzphlMY6oJO0e2zn9j3eASGyJr7MaL1hj
MpbBXe5D64Bt/EcExx7mGADaH+P4Lu6c+WfF3MnhPW2TtPOwsMCLoF1TvXoYiZ86
B6cxXiR+EsdoW94LHsNosPHYQRv3hTSzQ8BhVqtuyiqDUx24c7Vq+EtoJDY8xEFf
BeFTpcT+SL/a9swXwqHzKBMs9b/FFgYIG7u9/Y/ruZ9KpeV7+84NsU1EeZGip83o
gctAm7UmoM8r6tF0k80hiyl60xLkrD4lYD3AZUQSvqyz8qHvp2vcQzPxUFRl/PRP
y1OJw1sDfBrsvs5Zugr2hpW/KdTszCmSRMlHKNVU0PHHGNaIPRJ3w/NMQ0XpIV86
2dr8sOECEc3RQUGdzCTdiVi+l7rlIj+RH0m6usaPM2UhrcOb387wZvNKpJAI12Qq
v4pJR1C7AS2SSIM3qTSMEpAF46DXEodQeUX6LWjBI7Qxsh5FwlI73BsE9efyfg9r
7otgSj1PuD12VX5z5dF4+bmbycnkzo87cOxce+pknZ9aUopeBCOMhDrynMt/M4jb
WjitVMt5J7Kr0gyMHjBCqM9exVWgWYfazWFj7Sv+hLutiDB02u0hUMGbiqV3RzYk
bsbw+uYEkr0QUsyR4krxH73/k+YOBQXYDqdy7fePNXVn28Cs4lhKAwOeQs436ExX
Itiwj97PNSgqaLWSwduJitytV6gFBB5K/UuJjnmHKhLMGxJEeOmnYgLvMaPbgKfK
d/s9Q6Xl6R1NTKkYX30z5Ro9LzGyw/rWPEpfXeNkxD4QbBvaW+PUocqeSNfr2nLJ
1KiJPynsmgKKXjn2uYGN/XNj+XcTTx0bHyALYMl3G9zLnUR0hu76nW3lwwIsHki4
6Dp3QTbnphmv41fjTBr/m9RVlDuTIsAGEN54+94oSPMeD/Ml4cN9o6u4tAB64qNn
xNAx6RJfuUmWE4+ctj3tHWDGlJAxsrPm8eNJ7XoPYBT2Rks67h+OgCm7L9F8kTKZ
V/DYaIaScpiNBblNNSQrWC/9oloRnc5WN0BgMbBth4oYqaLWoK2SC7qqj/jTShor
b7x4s+dXSH4y6GM7n2tfyvbOYX52jlLUhtWlz+cG/Vo84NJfurSv4wJ0uguJgVTn
XCLPohEEd9E8wzSGgxSpPqDghYw/bP46WHA35+oSJShUVjsqBuvZVNVsVa7cnqe7
DVzd2ArHteKKq1OclenYI5obqF86TYAAV+2krtcHdpBrTOfDoXORzjzyAJ5J+t57
4imT/7TQj0dDS3tu1Cdwp0f6X3dfTQewG+zSxAO3/LgMj2Uv95AzS4Lq8rxsc6ha
9oxfHbE5BpoOGDIO095D65FhKqZS6rnJW+4vvMY70O6q/oatOGwNnxWW6Fbh55HP
ya8A7gUsbVN9cJ0ZgznfJEqSXsBFAIqdmobsFRSrDH4T9I42/uhNvkv5z0NUP3CE
O6h+YHBk29XaRn9M2kWpPKrTmgDI0OUp31SbwDdFIcC6wFdLvphqkuPsFIN51PVM
Q/UUKmmyGW4swV2HtVUURYk+0D6k6JT3evcaNV7d8B11rtfL6ptRfbMcalKZPwVB
6n7dDMSUcfTMLX/T16d1Bjj6Z9bD3mYE20OEn5Ko+tPW6vxnlws36BV8DcFHN3Im
ewcUTCMhvnSIkeFrZpvvOI8b+wCay5pSyYa7Iq1vB3C+mN7E6Fi2g1wqlS3cdF8A
QP8Z4iN7IzvDWwellKEs11q3xDDOPHQy3Rzxce6A1uoWARSxHjLNxregFRNiNHba
UNFiIFvB4UTPQxncR4muapErvptH370knwdJ8AF+NWBpTNYxqdNMtbTGEjQLHGMO
95UsaMWPL7W5MfpBHAGSlhUTSqSP9rhYXUupx8DMEFCHLX4ObeWq1/lY4xKnLYZJ
wvHtJm/ZLqNnRSKQn3fLRwI7Bs0ZS5VsnwBi1XjjMJX7jqx9Ic6KnBT7To6ZnEn0
ZAVzt7NdqstaEMkcarLXuEJLsf6Q2jIqzu5oCs0axAFVt1AYSYqt6UtBE/p9LjWJ
vVjaV2P773+s+3U0QxPlNeNY4hGemyXD4j+NpiZhMnWKZaQRdegvGYPxWBWz/JfS
f8mcYN+2WFP/e/dcRZotqF5mcxHTQy//n6pPsyIuCrUAb6wEovF1bJeHLJzopeAs
ta+V8K6CGCboLs2i4NPigZBDFlCKAjKPWboEj4IouU2bEPzSb8P2AMCyNeywXBct
bqSRWty9i3ltcpvgi5ZiR58/wn0U+izhv/LWFnn61QORA6+KH3dlu1SxyB/5tlWQ
d0ggpH0zD7UaeOjwN0XKQFY/Qm2U7y2NMTu5/R8zCOwiaiiE4rFh/ogfeLd1paUD
p/9IHSh1WpNPqWAQUpLrUQV6uAHPRawIMG5LpnGfg4XEtPVq5CO4z+SzIo6xFWLV
DtjOoOYlOBklis8y1vn2nmZ6UWE0VQwV2mR0Bp3i9gZJXY4ylfJ4yhfPmcKVzrOp
xb25HSDrKhsaRYE+Mrwq6e8Gr8CzMVSTLpuzCBn3f2477qzOM7SrPX5njuiJ7J7Z
G3a+Jqt7MvlEeoVpcUJXMDM6PWxiFefOY56T8xQbfZrDj6c3PJqpRdsay7Ep841M
LQyEO4j/4QQvpf1F2I6//v426i42dZyVeiJyU6CFAXqn7nKeNv/IEvgenkPnWaEf
GwyFCF5NTYDaiPW4xuuMIHNytVaeo1MJLneBBreUtwiz0rYeeCazBsvwPb7HRfgy
NDD/VIiO6Paa6uUjfmsEjsMuzoO0wbjfl5nVu7sDhwuazURQjj4J8rX7xB9WNawr
oLuUedAlPSYQ4aX4A/NoY93VO7MbTGZ3rK1Yehm6ebb2HOs3WjtyfifXtebqH4N1
elzehPlQHNjthCcs+hFJ3Y7cYj5IaS3IqT4jdYvRxrmi8PkvedIAV9IoPVkYabLc
9qlgpnPR7GyZAR++OB9xmTwc+mKp/mlQiukDg5wgTsCPB6+cwStcQZR+j6Y3aOiY
sz05y8O4wc/T1yjvTDeYzG9ZT4XemlftJYV6DK41CZs7Nfsj6SJdJ9BuC7IpYJuk
jXaZAQQCJAJ0JHu64VWF4vvjl4mTmAIwe8TQ0NQfurnkDF+7Hs+32/EbEm1I4bkj
GlTMForR5/DsbU0CkElZzX9ozCHYiHKS/kYPxyfFYTSXekiu+4aNSjqjhLibcnG5
F4rzLmFiYtjac4g1vNTVArmEjxZkkFzwPuVj26stVo+ubX2PRFjoY1kqdNEwaOGS
+fRuLMTBnIWs9l+i/0HKnvXja8aSBhvcTto9H+pyoBazSNexuSQ2XnOJoaXQ3aNO
hB6b5ECSLSJVWkCikf2pB9ZobijeB2dCQ+/digxOSekL3nWDs8EdYHKjau7qD377
dY5h+hn9UYdzWpMOfw0COpP71ZbJcktWp3RbYf0xPbYGRjLiaxKVSvWZuaX/kgEP
4nh2ym8TEISapSaJUv8V5SHGr/0h9smvubZ1dFdnJHuFg9zVdtxK/Z4BVRxcsiOG
xRUsDAm8ovS9b7nIVTyus4e0S0xb8Ixda1GGczWcVeT7Tgp57zq+6G6z/wVzreUN
mTi42fijNVEyaO1Cdn/T/XKHhqJl43LIOQ4posmDs2Kq5MmJxaoEHo2TFGomPtnC
Tni/HpcPtYV4eODp1/UnFIDCJLTUlxOOnMWx+fDA4Pd+EH78jt8E4eV0e4qmDZ5K
0gwvWDd0sHBkdsxUkXBO6py3lRmx1CGBobC4hDo4pLsfBTM5NKZCLYGg284Az430
/0m6zmamLlt5nzZC9kx3/FBnmuh2aUa5FrRS7srORA6T9kzJfPZr+TEpP4i/KkKA
HP20WesrPpwVF2zgAM0SfI2yD4+Zh9mOZbEHEAbI1XRNGwhqoyuj/e75DKN8a16N
mm2zVNuZaCUZ860j8uJ3YYfropbZ3J/SeKCvA/slFTyvsYPjlauMYEfbKv9f2axd
84R7H6LsF+FCyorqRjnRbKQxBxJEaI2Gi95li0lQu4DnnP+MrtIGMSy97Xw8YuWO
lxOC0X/ZpLIpHFls8cbdwyzZCCivgA+NQ2aVFLRDGhhkx882neZSunHYi2QgLjt9
rgRg1ty6NBNX8PWqdW3m8YK9Uv+W1NPSi626OQ2rar5EO8o0eL4EA6v0DlGnm7v3
ln3mMkOplTEKV8SQqmWZl/jsuLjPcozScN/EFdkhQPxNGCsiOH1uhNmqJF7YjVs0
bcNq63u0cmU4pWxacva/Z+Rvb3v+aV3VPjp5UPouzu1b0gKEzrDSnyXbs5aYWS3I
J0/zG5U5aa//Il42nondtXVkZ1TsSlOWrmyveaCglQELeGb4+B1tOGCLSEUBvGWm
uQaLaGq1lZw2xlBU371BXkdxsKnOzLKqAmfw53XS3LIHJYO+CZPasurXAfGYF/lU
fx2Mafp5A1O91ex8mOfdhaan1320Kxl23I9xp/V7NFmKf5LhYXtmsrG56YKkb8qi
FL5Ci64KLoYfiRtbrxEWh60oTdc/hcxHfsV6xVlzPc/a9xovej9Zti21jJ4vB5gB
4GWuOezjbr/KmPM4gFdXOS3K6jX5GZvtRe5jk4weKzTB109hP982XpbSBLuSz7cO
2s0Y9O1J7TuW4j9mNt99+iwqg6fX+32QvfqZRUvkKv8TpYRiG+Cc2f6FLmkPrRLA
`pragma protect end_protected
