// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:00 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pKAAfmRd9JyhaHbKLGrJYY7dzrfy7QByzJYQGYdK8Wv4qDU7USGUdOLR2to7qTbX
7pMHGJPmw/F2DtmizECgLIKSC3+uafGRmqS2V91IXhYDAPHGj2Iuq+SQUUU1qnHA
ltw8razZCl1xInTjrh9A6ayALBViQ0oIh5cp2/tJj0A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11312)
qUO2PdYjt2X8iw5dC2uIviNhZG37ft9lAjh5DmEfDt8K3NrP4SQsIHJReKu44BwU
Vfnks6f82PLy4OQx3r/cLso3ROptkuzduA0NknLgqVptoqvtDNTLgn7/OwHE0zgA
CPGgASu5qnWooEFMhDubIEGLDc4e9GsNILhL5cvqNTzkJAs68jWQzpzglq3AdScd
xA+D4j4pS3enfDfYD7Rp8ImVBIM78R/BmXSXG6ITxs/QaiG8od75HCGRdPPEJt0D
0s6qiKo0CvI54r7LyrzEcViM3RyDCb6hWcFneUgnFp8T+unmgrL7wFFII9QYTycV
eyYkeRWuwB8+eXBHn5UA5Kxv4pzf5QbuaqhGd0ly/U6KplA1xXvlvtR+DZAamtwD
9EzKkfoJvK/fyaEmH69hMhwrAwL9C+uqjkMawKMnM8y5pKBJAsDr4KcsXthDPE8m
yzXAUk3g3jteEf/tcj9WSKkpF3hjzx0bjLX6BpmGSyhvUriGA3bZ1Yi69EOndEj5
TueYhFTCL3G4PzXaQxo5C/9ivtbT8BVGv0iutDcOpYfX0X0njgJ8S1TkVGmPm11F
XAjH0BTPtG2NsRG2wL/Ik6yYjCxaHv+aGlCa0XoyeNcC0hiHzWvkuIdrSVKOHWaF
Qoj0GJ/2fclveg60Nk5vfcOHYjlKzmgai4V2CZXe173gYsL7lXUoy+lxb52TVxRl
2IWR7NAN76NDy2CSrvJNSVk7agb4OzMo1JTIPMcx//qmHS0ZcbfoU9bMpLW5qAj6
5B/E2cc0NCLv5LG9pLE3ifT59mvafhCsICDErqXwJplGW7t2+tctjDXPbWx7usxF
3H4DJdSVkU07RVCpi1NlrjCunGJeektAL0IrKmw28ep2BTJOMAl8XC/H9oSUaf6C
QrmROYV6N36TZMMMRGczPkXveS5+vcI53VjLzvEnP963d5ZAX+u+op2qL193i7/P
o7DZImk+7RJ2nz97cWnJzifhdeiyWSPqHRgTEo/fi32ocxRsyp9bo9O6AeVVQaZq
DDMRtCtt8V6h9QnshonrbA1RZHzqKWsb962T61YfSipTX1bkhFodAtw8ZAFOh4+n
aXZUARjc2BUvCBfG4AKZcFItqvecRBF+a0RZNBAkmi3P8MLsoiZRphtxJTgP4lt+
VPT+w3ZjzK13F0qjUO/sseZ8MX99ABrAN4HPXKvlcAMzkjPfvQMc95i+b+uWN+Y6
LE1bP5uXK3dRjBWEFRx/u4z5mBZDppwm7e8Usjo42FyKRi1DeQdZYpSsGTMTmLZR
oFdMtIHWQZNj0a8k03wTWmP0pBz++jyMHHvuIRrUWcFHvVgAaZ87z2DTO0VFVp+s
p0Gvn0TyOM88taTDcCYjMi9uHwl8H2cAcj+oHWOannJ23af+X7kVIvqbtanxE4et
Zs9MsB41IGapeAqaRaqJrWnl2zVcmNTrVs8zhYjbRQvbMbAIOAK/8ts1caMO3ikI
5Og6l2iSSRRnKMpHRz+3nW7btjUCW9vFEybih9PUUMz4u9SPppxsdHXu46fOWJVW
mmawH0T7D4vYapWXl1Hwsjc20AUtD+/xzz4W66Q6Z2VKjSPdkC20VZXxcYGTQugA
LGoxfqbgY33gL+zWqkZEnvlJBxo3gwiqVkrKCxyhQ4gkP1YprgveUqaLTHESiQUS
N6lxsmht/gbrxgzCIue8duC6d2jiVY1Ufa1dHyWLDkKsWeHMqq+HONUtKmAWD21x
BNJ87ee2ewFeP03C6M8hBmRv40EnJdtqvz8r5iXBFc8fESm1EO4xMxErkm0htemy
Rb1HCeqluutGEKlrR1hCQouGdMB5WFpL1SX7oEuWVI+v9ZPvvC8YyL2jrXoAA2rU
E/4+HeT9hb3s6oXDuSSRa56w/vMtjh/i3YQh9cVJ9+Lnj/GorATGUnMmOwqwHYQg
h+IT+maLktU2d2nK6HEyBJMii6rr57hlj3lElj/UtqV8hvAcQWGjsA94mKAhymY4
ULLghlEKaoKjtYRWgyOCF82UcfYrMPOGWwHkIRhX57am137PfiBW5WMLZ+8JLREk
Wy9PqS8QqoIHxQI8xXnP2WFLTg6GbEC6LJgzSBgulZuxTwhmYcbwNRT0bE/+6Yfw
nx4M4Zd6o+5Csl19YOMdhjmnEnoDcl/nwQGbunk6Czl5bA9zdxlzzL40wLLC5NQ4
XjL5/SKRIXxphXgudyhWWNc0TIVv3GFw0T++yT9HKYvGzQ2K9J+fFhx3PxSYnd4h
amCrXyKt9FeIRXJwGKEMRu4eh6tOxn2lQkh4bJrooHpRAtwGPqtEQJp/nO486f7f
aGVQUjyuEFGEOJtFdpdpeXLZ72UteNzkZSNEMPvRzPDeycvaf39HSjUKvtp5lr0L
iN73oHlLZns6hUqnEtghknFPKMFxjDbc4F5i6tlN9ZLu7513GQfuYqECIILATnp+
tQzl/UoeB5TenXP1U9lyWaX6fuv7Q36wKO4B/dXlkIjNqzFoe5HaigSawJD64uIW
IYkSnslmP/igZeeV9ivNeFLvJ9K2I3Sn3+PrrMXMzIZ7pg//vQfoN4ZW6XRN1SJJ
Z9rxOSlcV/cL0YxyKqc1ciEPbkYoTjPz1+IxxE9QHGr5yFmV8YHhskd2mT0FR83U
0WGeOcjETkKEYkS6XhArx5FRaigE7ta6dRi+14a9TwcFEeqsaYxXtDXs9xR9mg5f
NbbsSOE1yj/vUhjwJ0uIMLdMfMLQO3xsglk+jV0mAkhvpSV9fcSHvze3zirB/7bB
kIxEmMBqU1mdKi36Hthkg1/cSh1dZa3JtTWLC/u4RrxNfILY80acGVT9TQ07TaRQ
fRqYwz6ToixisEkxaUc20T78Vt4TiIDaIbEZm699zvqTOHhu6uOMfYVp9MHPp+QW
+ek6ct++UpFZFGhFGdykm5f6n+CjBZ2X4fLPDVi0ory4/pOOf3mPGcRII2HOyC6O
NThcNHbhYBdZJQeLQnfWi0UbtorPM/UX1UcMl1jNo+PhVtYqMNfsHt0bfy43i1TD
yRfCtofu2bnliDF4oqMW26HI1eQqZZACx9Q/r0zVPwsYLTHN7uCi4bFDQo8QysrB
VjxxBp8RlqaQa3gjuDaDuVxLFOQ+8XtsJPFWsZrS7aSLY2II4Tpn5IJxupfR7Hmm
p+sCE0p9/V9LM18BcXlI95X0DJa798qHY1RU6HbshEzQ/I2NPY23WTObwT1GbHzk
UpiZtImDHye7Lc4VwU8fgwLB5XirbtJyJy41MZScj3sNZlYAihxvUoUPYgqei7t8
4Y9OlIO5gzSCg1xyRk4Od7pLm8k8UNC8rxfGsl0bMVslhvt6NNkcBl7MJ8AKhIKq
FM0oEWT9Q6cUqm/xu2foKI1QHI8Beohz7axmC6o23/d2CmQ2mxz+xPTiLSvzxJMM
5wgebvuMrHYwgtt91GStfIz97QfPxtAbT2aKmfbn4T37c/vg98SwNVWtbsWQ1Hkf
2fIU/olXpTxArhoXw9BKsBByzI3BKHlyDJkkfWqilRzdWRL6vMbl8E0buU6xiHkk
iGlUPwhUL21exM1VcwRMp4YCdeP5ySMg1owd9L2Lp26asNkPNl2zENrYm/8pRLGp
LqzFKYhQSuiEuBS9rU5ENg21bS2me7ciflLmq9eedYKSfXsRO7XLemuVXzrTEOtj
BG/8BSubexgdLXJUwl78IHQnM5jJAhsTsJIpyQ3iV50d/RSKrzEPyLGvG0ktwn4q
ugMosEp48Sbp9whOz6+klbRXcHie/o3nIvE89x83L01PUMza1VY8L+tiicZ13tfo
prnpwvhjcjHu8d4gTEaN5Ih99rlMkCf0D0wFIFai6lp8WoijjnqoOpiWrQdd6KDN
KlZa1V8GDxPabFpdf21PkJiwz2J0VZq9BGGZguRqhVb24EWV+0OlzvomMxB1u0Bn
Lrfl6Z1MFaNgyhP2YWeEn6aISvZ4iKlntxA3uGIsgg1pu9l3pMI7zdTq9IfbT24G
cHwSa10fDVSVEPzaMpM7+D3zgv2eAtkotU43F96N5zNwSvNlyu6fnUMuFqChd51d
d9ubFV5FvAnOQz+bTm7yJJaxFrwE6hYF/4F7URfoZWPdcgyg11fkVwu/HdjDGh+G
DMwT+IZ2uKGZqvaxUfUXN6pfGkSd+IPcWYG12lcv2V02//m1NSNvLpr93Hzhj1Fh
ykZRa+qV9VrpMnX6TuXfp50sxnEO1fKDahil4jA1cb+gGJx313bfXFfI9iqzVdcb
RCmFYixld4K/nZMbdK7ijpcplUh+hv+IqqQf3JQDTSilAZp1p8R5NnRDQyueUEW5
9Df+pQRLJgND94aN1pmoYtEvhN7ssm35LFwZMPsWFcQGOET4jq2OHe60d4NcQEZn
ykUrJCH8La5UexDKPNavhmGd6mdT2b+liXG7zgFDUAHJatfFOGmsKqOT8//+NdPh
T+p+Rgwr9JExPQVLAzqjXgc57z4vFpMaxIQU7q4vnZu5dAl5sxcRvabVsPjG0o3l
thNuXXm0EeLiiNAgee84EIGTGoTBpyT7PbqbOloC6scx86ee0qjoiF+mZ5BmOW3Q
G/PZSTeTnTuz80S/T/YY8Tdet5DuXJutkWIZIhC4lCZvbjLWOzRTRyq9jffSF9qn
K7nd0+Tu8y7TwFBep9SduJiJy4/2VJEaxlorSQmeGDGLRXhKJW52lcXVBSCFWxFv
FbMlQ+Wg0PebExUQ0aVCS/oVr2X3g5EMS+lvwkTm8eecD70xZmDdzx0LTUFGk+vY
ZcL0lgGwv+uiAiywq6gwC8BDDGGYCxhNPvwuXTcgsuIgu1/2etCSAjJ/0k4UR9jI
3NtcAZYvs61w9N0+tNTZ+tTqMPPkqomWD+kBIBHdGcxizVzjQ8A7q6nM+tyTyxRs
HQkFWC9QAWXTAkzSPN/o+fWxuV7OQnCjDPkyMjtJwPPg6xZnRNS7OmBWDBMnu/mO
8YOKD4U7xhTljQMN9G22Ce3ThvvwixJNz9EQwUEW2qqKSEt+CEVp9foeVIHFFE8u
+3Ug3Vci2MnObXDFt1wEe5pU2sPPSVWj6vFdXn3qFbFYQo9r3Pfg0gtWyDpsezNg
cQYNXusPOZMVve4bIRIs9cRUt7n7AkonFHzwB0TVJHXGRSvEtLTMOLVUaaK6S/mv
M4dvW4utDloLKk8wwCyDXbvkTdq3cV56nChwGJQtijdNAZQmjCc7CyUC8eBEwrFf
sxIN8mR4mGq1V4uTk/t0hXKaNq2CFxW5QecIq0DlMMI97Tx1zAtOexo1Qs8HlVMK
6JAY/rV4zow+aSoDlMA7p9d5IgklUl8a6P2Kz2hNQBo/u3MSzYhWHiboC/5zHQ4Q
HIOWU9Tqy70ufPRLi7I8uTijtNvdIhSQgIuEA3N9UyfdmEjbIe8ec+f88rZ2eLbe
AlSepxDyu7Mo2nR4QtDc39BVJLqESN876JZmj1ZpB8lRgV9V7NlByYmLLotbQTAS
OdSEBuKD7K+gk0xdC5uryN1hltncqwnJlcrdyCSyMpt7BwK8cs7/W5u40lHZTH9/
76DnSQKmpW7OhB39mXQ9BBqN+c9sAs2MWK8BqCSEedu1xf5KRdD4by2qV52z9w7F
8vpAYhOsTouVjm4fLaQ40KB+lLlfBlVacCmxyvxv7JJZLU66Nw1sLj+UYSI80AOP
SBSQ3bE71nxfcLKCVW15RnsFk+hDiwnBlSVk/162pSetDGdoPtWEuHSKdWxN0H4E
QJ31INPHxma2akHStvUEa8gLuqb5c7JR0lHEnzmFd/gXp5sQ+B212IP/8lz00WeY
0Lms4YnmWKyfX1M3TFac51CibGqJ74WSNp1Jpr9bAq5z60pebkVlvq7j6MWLEcPk
p+535lxUGDEJvazWDMRgFqm5IA5PGzLH7UW1sNb6N+xloOlCZ0C2qrZT9Q3ZAI5f
LHYc0IC6DwdkuNUBDyKk+TcoUZCj9M2kkbSNRR33THvDuGJw0bd6NXC5xoXq0ttV
6HjS5TvWMWBlyagS8QgSWemn/4HA7Q+lTlFqU6fEOYd6YSQbhgjgi7qLgSN1ddYR
pi85xv83gqD4lRQ0Utf2B9T1cKxmyhBCoEvdaPRRT1f7mGpkcoVREhcNi6FZFbiI
xAco/C42oNgQes45RXOnqGS3oSoSxWO/yjt3ZmyLVyCysnikPsDPAj1548JsT+Ds
lXiaGJg8d8WtisuQZ5S5A68FJgJpkwA9hKbYHPMpF58JUvAlkdC/pc+mtYNqI47A
VG0+RlyW/4Vc8rB2wJj3ck2T5dqFtfbTcq24/rzpx5SRK0Fn5YBRdz6NJREf7m+B
XqiAT7Pys9iBCu1EUJ4P3Pj0RXgX9wLcRv9s+fFM1qLvznjZ67lG5wRfC4u6M/Dw
BImBAfN1OwtHdGSKQtjc5o9yIRcd2hDomjViPWCkSEe8ppAFSRonPwxewmr1Y09h
UGKQ/lnpOpKMMBNbTCPeXp8xrFESr6+gj8Y1WW1es9Y2bTrjLDE+wYmChSQFB4JT
H3oXQnsqebAb1bHy0OElJs8C+7pc8TMyi7zkkXFULYsUC5voBtft7jX5vMKZZpVj
javv2WHeOqeFCMuEBTI65TPYmrE2HaoQ8qKR460iwzU//0FAe3u9X8NTBgPSrS3h
YiPEW61Iq/ELEBrPUnd6gCX8kpXzjI0YxmVfnfd97QVQzSpZff/vg2vM9eRudtwl
dnzHUVhuF7h7vBwj7YXzW4az/uzGSQbVpYwroZW0JjZwf/pr6bVq4wZ646ti3kwU
sZXKlHN98IlEj3zEcV0BJrQkzWi0pO471EU8ZQlzLZlzlkZbRN5abXLnKzSSJI5/
FCHPUkjo5SZvfJYdJ4m7vSLPjTKnmEbJhvkW8UiMfGYyTcnvRb4bbkBlNr/6MgyX
+iZ35GVAJBt8Zoy29Csi6OT0lpJE94NGMXSQQYiIFmnSehZ27HAja63AXqOq4lVb
iGny7wHMKGh+j92JoNzKID14wCzJj5p9eH9/t8P4uj403MBZHxXwkEICbiXstG6Y
zEph1DfchyyjqLig2WSIXZDQPKHdju0BD7pivIzj3tkHXzRNkfsUKlKAbYkRtBQ7
XsFkusBqOChE71dKVgm61jS5hF7Ga5zw1dlFpl72UWPfRDUWiLfcEgfPkm655Oom
HaXlhpjmgVV38PRBmwPQcQQPgtOhpcMKFx5FbK4510p9iYonAY6+XjnpLHhUvUao
A7k3beJLigrDSF7Fh/Vv9xT3hM4OIqXMu3Pv5b/og9s/OAkHgnCutxL9l/+OrhW+
XK+o/t0KBfo36+BpEhU3Z291tT/HNKr4oagWoWY+QqZI+pEbi3Mp4Xs/OP9UQk8A
YmrG+kyqHWFaVX+NlBmN2XPY0TPNKM4ifsXtiUGEqhDoZ5vu229nhQjI3YPaP3v3
Lf6JT455WeArClHIN4xTchlUIjZIDifq6qaxwGWtn3Lv8cNNMnvoO1zpiWNIS9fo
g/807YA5oCazWnOOeTBd5ZwqgYgzfbit7LrZihJ4dBGP2NE4ZA70VoXFmKgl5EDR
FP3tECiXExtyHPUElus5ZbZ56z5aiFBnYCQ/6TQawBxOLF3UFfB/fZBmYBnjNb6R
fjukChsF5p5ZSG27mAz92JdPdrh0yaLllPDuKQdByURHMlEAK4JFNsUQDayLnrQM
yZC2DDktbAd4cf6+8+ULpR2og2/pwS2y1EQR9oQdxHf4TKbiI5rkUgVo9fQxZtg7
TukOnGgmrYezrBQfvsPOrRrxAD23BKOaTb4j6PNJKyy3yZrWftkrZLf92S7fT7ya
qfbfHXULcsIimK//bTUt9J2I23PCF/tEYJOF6nchJeCEUc2FO4f5O2sBu0t0JWo+
2hrQ1GPkZ5Qz9+cwi2FbD5USTd5g+KNvnZ7JlbB3WrVqJoeN02H4QHdGPc1vcO4c
stI84d9HmcrsbDQ787GuAEwiEecUplaf1kxHbbIBS8xghl+VBiZI4sUeDOzvQUJa
x43hqtIe6rpweyyA235zuwZJ0Gy29b2goEvE1ZITWKypOiklwbPh6F7dB5kyR3do
mkOatahPJHA6aBkVziLDfgMhjIMCHkMfBuYAaea/LlA6SGvGkqy3zydxya1OyLli
WgF1+Huq0/dde5bY3/y40kwFTcI2VzaGVJIZJzf/obcQg00+3Abk4YKTGZgaLzdM
7jhEdoqUd3yPaMZK06OgBLkDorG3Q/RLfiVosW0BFrTXE+Z7IDPIiivfcRqZ8Jl4
OjWhyCaVpdt9HIRyA6u61Q7DE/o/Zk3SwNUD+ew+cJcfmRXGvW6UPMmlEzN2cLgb
JD2drkxqGN6TiYkmtPgbxe5iTit4CcwOD3M27Gr4jCAsNbmE20MmiOe2MmF7ND79
3a+o4OeApPofct5fAxXuOn6YsMe7m7GByLCppxa2LwUBCMR5gK9JAKZ9qs6l4Cgi
ES0LMBTf9szbCeMfXkY2j5jVAPSqEVp2qQFCHnKR95QKEb4Tk5uaSC/1sOZCJ+lZ
qlyCndqubFK9Vp7Evw/VkYzADTXByupOJmT3CX72kJVxW9QrAGtAeaE582c/5qpq
0Nq/3c2kapmtrOuj3xXbPyw/H/b7HU6JHOa/igVv8q13/JHVqxJO/WE2mVK3QtaG
CtqMHdOrSqxncLLVweoiVafJJZlwSTAQ7cmuJMK5x8A4LfQsMX+utQD92rBPzXPe
b4P4j3B0oAD5iXOlv/9gSF4fsJVFd/I60q0lkxGxCgie+rvE6dufpwLIMSBb32yo
oGt6X55ktUYYUIgU8e9aaE+dps3zDrDbz68lxidoE24KhHba7WCKZBjjge3DpBDD
bRp43zm06zLHjgNGwQsXJJD/ABXZfLnp31r2WDj8iZUMrHtWdd25QDmOgokU2KW3
pM/AN13jfjyt/REHBhePwXbwDzZgSbNq7DVIuYbSBkK0QSRo7hibRRrDHgJ9V0w/
SioF1CZz+ArdS2r8OH5iqorlZDn1ChYBWmIwRNaRjwnpSwveALcEwpn4MMdsUbh8
xnZ67jvVQSC++B2Het9MRQ08sRQ8LpVtBlzjmizu9Pl5xIXLUPTbvDUJzXw2DmGM
G7AWR/QvFs2q5F2VH47nrfzGl+GSJRf/isO8GaAFWInNSrWDh0NTe7tVTp1iQabU
IOu30Tk+4rfG9OkftXv8XSXAiugtlctgZLqRN4HxIlSIIXg7oxl4gtNTjZCl53wq
VzfCLOwyBpkk6CfwbSRuYabODKWUIgbpAsfHdeCDXkMtBxSBhtb9CIdxoXe7LjnM
RnAfb/MqI7kWr8wv5blrM7LdtOpn0Z38/o5dLZlkSEozTxKkFMqo7qZUeoIXt0lM
9xyFo40TG/2AmiWV65+rSoZnLq+U3st4IR7Kx10lGuM+TkOyDM3Tc7+l6ahS3KQu
5N5ALhZbn5qIPDNkJ039bjziUy4WqgKghfgxnQIturUqVYuag3VO6UbFyEgRKJQG
ZO2XpaoNJOTbEI+HLRPGDPhcXzuj6eaQQ24jQKLjcdXEROfU2IH4Rwe3OVCnEtHZ
MocrlCqAxWIoBD3XK+LflLV42c7xjAu1blRE5Hc1G4egQaX0S7YRNakQbw2a33Ew
x7oyJAo8phZ00MWNAbA2CqWnjbrrTF6dlxQQJzK/9VKUaN2sPjn8FkXGAJabsffl
uykOVL0vCB+07bdIvXpZAywmQ/L5g0cgdwvy1Q1shhDwvlOz8c+5MTTGTROtQHAm
BpfOyl9zGOzXNZhFZhaKC9cl03DQufiaMpb7JI/iPK/ehTULgp/viXGSZ4QzIJG9
MZZDWY+QpWZSa4inhRPed2WaFylobQr6+zjRb42q0r0BBSD0CBmquLX7iVR7/1UM
GTGNqR8y/a7HXk2SynkQ7fwKy06qVBVFG6866OsgXLgVbWAEm7VPjwMVcrPSW2VI
JnGaMEb/sG0RolWH4yDyPiHAHvtq9N3li9pMRyVfoaeCj3S4qC5E73dcqp90rlsC
0njUFJxt5TpoIs7jc/zHI7baArWH7OxVh4Nc3z7iqcOde9rfWOHqej2NMF8MkS5N
CRGOtvlg5k/8kNDiqNzQ1Wc+zzOROkPy075JK1W15g7Rdjd1LT9weIqv6d/KCy/f
FqDd154MsHrI9AU9x2yU45KXEDYg7LofR5SsiVLkwCExbVkb2r9hk71l6RczdnKT
q44fuJ/LtlHHu56JjELX8hMu7x7UQLDSoUBdb9QmKjDgCUz7HqCjXtUZhrNRjeif
A7g5cMfgpT0d4q/n9C6w6O/qMcqYoB89kpoB3m5PSGs6Q2qY/Bo+KhGazr+hppuE
bIxbkbrjLGyoNWBePKu0wTYv/eISBi4n/dSHKv1+zG18siNVaG3BXKmz39vI1hpl
x1n+nyXe3ugfFVuNwF4neReeo7g+VqjM8FWYYbOSi+axaiDPB1ucOSlJuN86xONJ
MupCpioWogvFh18l0WUAbJZs/+6eKTAsakWKgJp8CwO6aekk2F8MHGmpVrnsp6ik
gbsgmWl+DhPzVW4FJ1gn+Xzw6GQuaTSfq0dSwXGKb2Xl/oShJIWDRx1x28n8EGB8
sycJAkk/jM/WIaX4A05rXQT5LFGTP4H12fF58X2tzgvwqCyi4lLeW1pVsAhQ4aa4
067441c7OqfWC2Arvm/4um9FSIbgHPD6AzhMZW4zbmcnpWYdxeBm6p1kUVCs6P8u
HR9F77KmTalsbN/WDH6y4lv695JLRocCsCFIIS02IW/SSiuKumySDab1cMeuZ4w4
gl5GKb//pIekHr5A+sHuCoRrNZilKn88C0iiHAXj4h/51tDuY2bAgD6dNIwr0Cbz
i3WYuUf9Yx2K+M4JHpDZADMTIkzYlNAs4qzVhQDRdNa+VlNCTFy4GP1AsqTKdenD
VUdj1Jyj5Rl1dVfk/wz1Bv7hdgdP6PON+VcoJY54yEFbSYyapoLJgtV91DTdTxPD
qDH9+COxGhqqq9acUF/oFrgDvU1al99RtRS0mGa/BJHAtS+Gwh9lM/el3ngORseZ
tgxMr8Hae/T0YEpgQEREuQlnCZSdR+zGE8LFCPLcI6ysmAT4bpT/X1n5cPKJfzVW
RXI33CgXWHWqh89r1VnrNRI2wpxTF7qOy6Om4BjBSg+U+poZu320GR77TIV2DAY5
Rkiv7TwzoHfBJH2aTC7ueDBK3jZxsSuxy0GsUVuKBzChAQ0/fqJ+OUfs3QBjr30u
/WsO8Dh+R0zvGFYaq1YcpTdsZiQwbHN6mpLygk/+eofKFhVjjKUdT0vcHroJH+7q
DT445qZ991IqtPSbOAZkZDSN1oD8WBqFPZcjCSSBxYPJHqHYKsSFnxhQYsqyGle/
qCtMiPbj1R5kqKaVpkNA3ZuVs01tBG9PfRXIoV6J3ZKOQoRbmKvtJd3ECUjU7h7w
vq7bLG8UHHNLF7urfYFY3T8SjV9EhHKf2U974qSN7lxfhx4cBaoX3jcm4VXB+fj5
hXpREs/eR4rATMfAYbXkNR6r/41gJ5P5sGBlgjSyrAJmNkEMMliGpNSUsqOD60wo
5W99uc+IY3VxRwhE1AOQLDs341o5CnYUM2cYuGW+VykqqBNAdLqgYijHL9EainCX
PIGhiSR7N4oS4qi+n2hwTfv3eIqtV4KDz8q086BeBoZfv/6TuvriGs2lySl/DXpV
SE1kTio4FDjkI1rVqs9gbsJPpoKouUJ3gbgg9gqBOlFaDI6tZ1c3q2D7IbFDOBsE
nFHOH3quRovyDoJYK91MaziDsF8pbYf+4W/Xwbn30tLqy/AqG3pq3yFKLhx3pKy/
n0CuizTyqnpOhF4pcnzGHqN+euOz/L2jF73KsiSFFln+SHzL9ODNRSOU6gAdRbWZ
r8AiVeMPYmS6WpC6NtYZG4lhvbD9xDCu/qKfZsPCCXrKmLjq6IBgoGjDhbZGu0TK
Ececjhh/j8X+sDSTCDETqXwH+AzBLVGwaqOX9f0XcPcjCMzSi8VciRFODzdmNOLD
F2gRbrGnvxxl+X8sHMCaTqPEwBMC4BqqNsnh8Gf3tcU1hv9MAXRMyy3ehaviXB7D
tAglKM6JM32coKr9QCT0ddWBWI1AEhw1RHmgi5/id/gwgqtRJ03MNkZDMGDTqljF
gH6NsQ/n4MzOjkdCPvisaKWNFKTw9qZEjEwFZau+rE+Np903x5qCjgr+o1VzMrkn
bZaoDiZs6WZH9aDFMyXbaZd6wj2wUvh4WDJFa17L0UQJo1yirG7ukn7g9Jk5ivdH
vPrmpOawpZbRQVtUsgxc3GuOf85Lf3GRcfPgIiyTsCeb7lDKRMWHCv0nd7Wl7gJ8
BScwbCICvmF7mPuS7LWM+6qvb/p1RO5Mwqua7sojIXHBvRdAvmQLdMqpgZZvTsac
lFtk+Qn/khksLIAW+FU07EwUVqnEpkT7kOv5bi4Bx2kZgvS5LAeSqJJ/Iz5rADAk
Zz04YMkS1vHIeExchDbaJLfaBpaBRqDGLDapZ7OFeAwD+SwxYw684XtiFBNEYKYo
cOHyRJRmo/pcB4WT23hkj/JQL0nfEEtVMNVOiXP1r5mya7WZ4K6j6a5X93NhalvS
wOirlYlZtBjg/NaJmzc7GuaU/w0WtNMNI5PbQFvhh8i1a5r7IBQSlgPCMRPAaD2V
FZMLcU3pId4U6iJhDIJyuDi2AApweMd2WYOYzmzPbe0b8zGqpyGtZJFuswjNLM75
1QbiMh2tpOR32bMQVLCOH21WxJFOyIn+I3HwNK1fDnm+HwhshM1+oJ+q5A++Zpli
7jbXsULO9tO9SrpxAb9zMnhTBrC1P8YJG9XWcTXcCMlhakkjDQ9RFwAlR8l2/f3L
84Z6tKtDZaFc71jm5Q+MwIlSqovD6mC59bwE5aUxcQN6G6i4ZPv4UScFtL8+ydPb
YxDoURKGwFVz13XoombIDiencyG/HAvzhmcRJvb2PIBvxeV2FdfmeHSAuERddIEv
ABhu/ACiHFWEdD9kfRTYJFKYjFPqoTQM4Tg2R28PK3B00HVYXrhD14SfO46Jbd5l
BPO5ZABUgkifja/BZ0PB5NA8z2gJx+0xOnNPUiyTaQB4Dwf8EHYiQ7od190DpIqN
MpImCk8sm41p9CFno4rdveaW3U2Fv5/ej6y+BNHqIToWBaVnOehezO9IbRmQN0ut
6stQmWi5mGpd6RwsAH2+kdqYFS8ff7PIzNet8HhPFCym6/ZH60C+055eW4SAYghG
aIgjQ70lcbbYFCoEutYBd1wBIdZB6QegzlI8gLfWqd6tA8tDiFOf9KwZX4WWVWiP
0aKUnoOotbolf6xQPqaisa0hBgRm2rgqUcJxuR71paamys6fNGly5RbUxJPoBIbq
lhvliqammjqhziMd9zXyzQkDnEwLL3CSszUGCRQEWowqAOBvuaAXXJatZgfMtSib
phv/i2bJNfSIzvJbzVqW4bKK/wbcXtk56Yuf/O+cDFp4cSvL4vAI+P4+OYngPq8V
27zyldfhfH4K72LLGkbE75nVnCdvsry7HV9HIk9F4q28ydlV4OfghAMb2c9gijDG
os5kdUhEOVwQQhNuPpE0QeHuEzumgMcNA9ZL0bJjtGIrCX8gbvY2vCDmpgYH+GPX
SVU3ujKDanMOVe83EAaz0XFEayC/dt+mf2y7s6hToAw01Mes17okbIJWoHRt8x4y
Ll9Mi1JmLcv9ckpU4k/HPxx3byGwdARAky32mKkxpUMUZcQJkCpaGtlLpm6vQ35Y
W2dpphgcIvyEmDvgWKbnnx4/KKHKk7YHoGBU1WR7np2Jgz1mZ0qkV5QNQ/gpFkco
G+U4to/0hMN5UDSwxTOuurMq4pFA2LUW9OslCfwiZ7U/CUaYwsD7iZK+G0Wvc1zp
+7AzMk/T2CKnEFRW8VkQM8p7TGGuODLWmXZkfA3LjHdj4t7LlGYN66TWva9IHgCt
L+5xt/o/E+aeLzzYQ3db2WDeOgIs13MhmOx0ujBDEaWai8Zse1K0Uv06yJNDrOHf
eGejgAIMEd8jTapD1HRkSubnQCvn40VFCv4bKlySVVUZnlCzNfxSjqg6owThKEsq
wD2beVzr2Po4Xw5+lmuoXUSkVV38M0PrDaj9/82sPypctlP2N7bXe42m4HFa2618
EjvndqHFBiikUzAL8wqu0lFH3DVOkwnr31muugQ73/Rrk6rwXW4bochxgU9Fil4r
0sJY8jic56W97FDecCrIKIsnrQh1NKVGgGNPFOJ1dogEAycWGzVeIl6uUEWFpbDa
WYEO/VuMLvEe9M8ALgCi+KaMcrdYl3tV3Zt49wOmGfQSRX/iC/nlnKmg3aVCFFa6
Wjss4ETbujkcuaNMbWT4OigZHOjAbBM5i3HGuYlF/BtBSMScobDueZgDjN7SWJ8E
ms/SPNb/ZO812Q1iCmtcPthwRmhpAfTaa52gfVy5Cqfm6ryA3ctcqF8Yshvcp2vV
3Uwy+tNqtxEwiViqm5SCYLiX4JwYjEqz+lY/1FwQdYY/zclf6t2GY2dNnU63C9aE
Kz7yl15ROJYZaCN19kJRUy1rxXe1XxXaUzUnbYCuIKLSDoDeN2vTopGvXDDlQoKy
YPiwlxk513wUuzFicD6AmlMYiwpqazwfnw6lhEUanEhag4xFbilNhccXj6IM3JXM
C0o/wML77yLEd4c/zj/haZKDyvHhCqfX4cJunoKlduAuhX3asRFsMbO32xJrqryI
lOL+hCK+TLXuv2B8lQS5PW8bkDMT80KZbVeJBM2peZFKzGaDf2iLBF/WVWJDceUU
uBGMufhYZHCiJd9/Kozu8v4QofDy46ZKVnHuC0dQyH1DvjrBL/zCZVKKis6XQDba
s7oMCTKuunUz1bYHNF2y6VakJJSTShx4Np35+Cd8JhNBC/GsZHC33Hmx6Uox58Iy
GUx7xeUjnP6SuPD8dPVTOvMBYFfOJtWek0N3Q4cUxgBi87enGPaunlnM6RWT1QCk
d5EuGhWnBbbAH6aKF3Yx8BQCYlXG6SVPbQGuzWrPQsmztCV/hW+PKaf3EswcP8BU
RaDen8f/Q0ionKIK5FUi+uansY0WA0Y+TKXlY87T3eFLT3AQ91Q7SunAbAkNl5dy
mMvvDS6tLTNrDTQOo+Pe/pGReGYAk4m2bTizvb+62CJe/cXpPIUqsYhqBPU3j4Qv
wGad1edNvnXE94n7VwSp/g4y/KYpVPxWBnBoXvNiaBg=
`pragma protect end_protected
