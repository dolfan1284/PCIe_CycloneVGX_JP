// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:59 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KDmGeXRwz2u/IyJ/CpKBbKlyr+wIMkX8kH5dBcaS+QturNnlyUvG2lVVIDmU7wW9
33Fcgpg1pV/gsFSjw3ixMRjjuNYReANwqL2Pu/NR8cs/IvVQrnuSPTUOCVh2uKLs
ozszFGYuNObupw6Oe/dGq3egdYgyjhYfCrG00xZPF2M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13584)
i1NouZT5y0O0YTE9ix4JkUgxfAD+ZVTpkUB1XLP7CW6nneI20wXEzzcWdb07aPDy
cXPFJta7asHkcklXyoA73Qne+BYqWihL8hLsl2edK3eF8ume0xLR62X2LCXi3C3k
ULPeAxxZERmvunBgc6/ao60mqavXrirpUeqsus081u3rGbdHzNObGO8M10lOeP9/
4SvZxtzyUw2pXDSpoJBIQAkAbjV8Qg01gmePni9ebr4xVBvdSU3/oj9vof/vEZL3
cIZ0NIFXrpcA+JuokZAyai/t8mFkDGWcif/FI4ZgXYPh+CpA2JjLKY9HLMKV0V6I
iFwiNXyCZy+nta2EHgxBulEp0+/l5jkVspPjJUH1zaQsLRzdexVOPmBzvqv571/p
sJTT2hZWyPB5YipzYTKUMgeD82i3WA7HGbP1ZGKXLFYeyavnOOc0kFeED6KWwSu4
HNxhSxOAg25iDxVIVI506ZlMWYEcGtJZrX33bpz8SHIMUpHj3Whw4Tw4L4a+WCiI
OhQ6RRrmLPCikRkoofFhrl5r/BVAWQSNjQuQc0ZLfkOzh530EwGw5/e/7Dd23tbK
P9cr1yOiVD+H/x2PlWDpnYdeuBZdT3zDFtbVB9KU5D+Al6x0els4fEtdQLjVu8hR
tJPjcLYL0MkCymGyU3hj3rOtYGoD5WmST262iP89vA1cTlznFAxgUx7yjPQ7fN8p
yglNZfjwDqLsVilaL5ShLm85sdX81CAVWqbhuGxCgGWtxAKczBBIIbn48a0FD9Cn
/EBtfg/9UGiWtHGHw6MbLHNwUogldTIzi9Qk37JDqgVMDJDMwWlisUKQS4dPemgZ
+TZqFQxUqmlSluWFdvPuTPBtsp9paY8VbRmkMn+R0ZEf86rj4vmIL/tFIiSQTViA
6QbC44cMeFKgB0wBTQk0eb27aWYvAMUT5CAJfdTr1fhjXoNT8jUN3Xs8wZLM+iVO
Hc6AXzr0w6s1aLW/IGXJEVeu30Ee2PDrpZKHHjezA8w4lvsnzRfh8sDIOCwMz/Mv
ATFslXQAOE3wAeCggZ1Gb0YQ8a3Wlg4YEPAq+bqjszD/U4tt3y+RxF7QFIRZIeQc
eeSLOCIFMWRc/DVAtW3h/N1N5yu0g5WgB9Jpo/zsdldloWmwSQ9bWmZLd9sZ8EoH
skunEAgIvvfupvElpnVNzhvg2HDTnj1xN/geYe5G5uDnOEp/8YnQKruZ8mb6V8TB
TBP4+NERhNnB9vK6cCfq3Gw6YVqwMFE+4H5zTt98mkcbhaEuOd+Iu4l1ZXdIpJa7
nFksmCOxEL9LCeE6U8MxM6rMCWJEJtDXIeUiEOYfSCHcqknhzXBndMXACnH/S1E2
ZcTAKs7a1ep2IHdbMhbyqscRCL2PZNKhJa9aQw9ZsCbhq1IDGUOp1XiB74R8fcjE
7aoZRo/AvrZlC+S//gVssUXX1ApI2IoxAgnXOLdiPUJ70jjo9BhSZWr92NmY31Ck
4JJ8Ct8W8iF8E11k4/fL9pu+3aHSF7EYSwS29WoCZDzLPpz/jdo5TBBhIk6fYsXx
YmIL7Me0iZ0c1tpofAmtk6b5zsupqgGdCccRdUUevLHnlf5BI0frqOaqS0ZvgoVz
aKJz+4nyjHK/wgA78K2XTJJxzkbMwktoa+fuvO9FkiUxDVl0jQbdwh93kifkTkkl
5pN1Df5/oViqhwm9HwgO89rymrez/WT4XKrNbBr7JCoWsedNZa/1NUkz+k2R3VjJ
FtZF+mH1keCv/+izJAd+udQ2DlI3ORnu3MKzTFugEbrv7mTLIvhGE+ZnOl5EP6rM
nLRCMDvaCRTBphT/BHoXVV7Yu4sgi04YISI7xq4dDbgrnGMwyhrp9uunZPM/NL3k
FJITUwnn6Cyn42GQna5XcZQEycoor/rjk24PClsc2PtICyZusJ22pWxVXr9uu3jx
CpfMv+66azYg+oAY1K/4RO0azOXxXQInAJ15qctE6k+qfpZd+/mhjb2omFP13rwP
VPgGKP4akL1XFs5FyTbuELKiLk3RbOo5rvcJIOr70DQZAStigjyugHlcZtzmMYa2
97BQu4j5SS0/ZyNm4InxIUf2nJtDJ73NUgtia3qX1g5ydfndFXQ+4HA85bKmvbYZ
xDoeyaTb8yvovt+NzmwPyTKT0vwAfQsMquc/er2EOr9kVppyp8t3f9B7cqf99XJt
Z6obBalXOr3yg803e35p8K3/PTeDJ6eJ0vZOT/nWIUCdVND0E7FkVaVZpRVYdhMx
N9Bqglp8pNk5nSjLNh7dfIm2rdSjwBWUvmE6/wIZVf5+szSTHzTIw4ZrhjvOsMJU
o4PiAF2OisholF/nwpNEvmSj4MLaVT0l2dUTaZMniF3DcMH2g+GfjcKVMSbPCOth
AMzrbEW37nV4g8gtM9tSz3IUDhaIe/5lAT/s6yJZAwUM4HGP9myuPWqFLz7TqNd1
6x4ACT9DMRtdKo+sPEjFsZGBonUfbeWw9rsTOAVt5+0otoarQ5ac6Y2eEYN752qz
HoygwBqSWMJqeG4dYvj990XoGX7TNkavP3vLYhbVW5tHlGgY7t/4OjrkICGjiKby
Dj2oNZiCHR661aMYW1HhNdR2UU7P532bBzcpxGR5QU61rbMSya0L+NQoyZNi2nHa
xB2NMILcZe6BfrdVYC+BgfkQg3YGoOsge7zprqpxS3+eA8amwRAh9wyLqCicFQdi
RPFm42WdopSr3fGdJoEDJYLIz55ExHmvuI+16Q+xhDH7mKaaXlTEwwmRJUWkGCTq
HkMnWEojkDzHzXPOqDw/g9e3r7dSAo3wR9z0BeYnpbC6DmxPfBgKbcnhJGEpZvR8
Mrd3XeNC2ZQRRmFhATL3533Olf8VvgZ40g0vjN4XwB2J4h8/BokSjIx+kGsJKlbI
W6h6EnIbmbflB2kEPP/qwY9KhpPomha3rhhNc8ShyGoQ2AIANXm8lqD7CArnFyy1
6ShymS84WHgPEQXCF994Y5ozlEjEb0UpeWxjODnkmpqhAogs7yIpy3t9JXClCfSP
nfuonb4Jv7u7esXvegvmegqsqWlkhT0z5GBMk3z28ohk2MVWXn1SYaPe7Ro9endF
pp2dbU/lwRDvoLYmjIAzG2xo5zLT/eJGBdCpIYXaldpOEx6pL5/V2R7SBhQxPY2J
x8Ewe35kI1o4TtyplPTHTQSbJu2NP/7Nv1JQLY8gxGHZAn4oU2K766bj4VTEyTUZ
gLZgHZl2NVY39qcO9uBb94F3pCpYe4P58hHtsLYO3y7oltjAFFwf2YyfBmOM4PnJ
B5d/NlKqSdL9sxD3LnZ7XdKgRfwZs6raqPOTuPcW6iXN6aGZ91RO2zZ8sW5WkewR
4g3yiDapKXaBDT6QoQMg4rjclANcgmnXUghd1PwfHko2MtI+JhKP39OdOLIiuXnh
8GNbvSAuCY8tJuAhF6U8zlRjEk8mG1UImKrAeY8zmp9QDSicITyZPsQ/pUbaJtYw
PLYzrf0jh4CF0WY580VVm8U+v1DD35osGXcxrhDnRTwq+GF/M9/f4odTgEI3h0/C
gpsLIzKWrBwnKxlIVzGZe7Gqp2EULlpLFF8Ae2vjDFm5aIR5Ec8++8rJmRMzs1Io
oeuAO/DJqg68Tjg/xHarOHfDJvj/gxGBs5oWVS0N5I9rOnLXXusP4YxCHcFa79s8
SE5N+Lg6SF/6AqHBA6QZpa5r7AXqSUgP0OMbParyeQ/d146JVcLYYYCcQKsFaZN/
GZ/OmJUMPI7Ia8aTF04HHIYIsofrtK++/jpdpkjDxONXeWcTqXQggk3icYxRQ1ac
iJHWkSpW6/zmXF66kypGHWQYS5Vu24Z5vyR0eFqCHp+qUMCtAYhMjwwL7LK3LNrx
Zmad2G1kELZ/SAZcNCxxBaU62KLzI9UCmob8OJhi2I90p5kRapLgLjuFcS2Vy3rS
JGij4EAjQLoGNfkT7nel5Fy5FIEypLPE+ErkGahGxW3h0oT0app0qPcnb8xsQa4Z
wNdnQ7cTdtXeucw7E5o6cNaPQ8YFfkfFhfPlA/yFEgMH9pAonzPnQVnNAMCES0OZ
RQnMEgaZGDIsdkhWOcqkmGJJCyWpoCKyHnNiiYQA66cJgHX5BCuFR7cb8cL0Wmjm
AUQrxdOOaeTsoANczviimVKvNP6624UvzP3NDnamt65LYUE2jQO3rMgwoSSkkVll
Gq9MI6shkW1L837bdcBHrJzk0YuUUODQ1jLItXEpo9I2Rx7Bcvl7W1nFx/4jSWu3
vLliUo3Jb9BwG68slP38iMLX/cty58AXwsADLegb56iAOWDpZZZjGAAaXj5rI979
EQ5ELtQgPNHaMbBwcaZ33Kh2eoAG88clddpVS13jbgk3GKjGNW6Ki1kp1GwPKjxB
pFfOHNwLBLZCoAPet2VUYbQ/QBplVrOymAD+7uY3QKsFh5gAtG6XIccd60YXJvtX
o35MbRwXuKZF9c4CrquEurZ7/QiPKbBfiGblCRa8Y5d1WgU77V+8QSIOk4G/s/PN
KqU00iG7VqtgxxMWB9c1l+iYt4aV4fUsakeEzd0k1L1DTwmDiMyi+1ji5n5mPYzx
Yzh6PWlL302Df2s+TFnN5s49Bh052QS7TdzT/3ZspRfO6kmxMFsgs13KE3e/yuH6
3zQ/9kbrGjDIhzz573CSxCMV5CT3IBRSWpDFze4NxrAtZlswUgnkyvf7WsFZADfm
7MPA48gwIXcVkTznXXQBQgn9aBv/x88vSkmhYw1KMgk/Ak78QNfgfjgGSSN6NkrL
vvD5FtFckJCCw65NY7iR2w5HgEax7yarS4Ru7Ragg93/0YAr+jtdDRWVWGE58P/G
OB0LZMfP1rs1utFkvsUvSqDo8l91qHjY84cF6MAM/A7TAcBM9VRPus4zPXS7SYXB
66pnSjPLs50m/ti+sS3xcNw6+vhnKighYPQSsLe2d1p1V/iteyR+KdwfUaKxLvSu
+CkRzDYFBsvcPKrrclwh3JKMZztvr5qRuLjmHvnNeEvZxvyCAQYHeaVRpzaTEk4Y
6/sgj3p5z1sevetE+z5Jfs7w9xnDG0fVfnDxkMkeaBn/Sr/zap0Fm0zbNUPe9IpS
RT5mtN6LmRdUA/fwRpjzN7+1RmIqzXYpwzyh66g/2bheRrPdewNE/fxlGEE3DTeP
91ezjDszErTcVUjPxCoCti9wOiiR5dBDHfZWpiggFJ31zwInizm/2kosvKOlJGx0
/mOLDAzuAAMAOgWDTbnWg+N1x1qAGoannMl3SkxbbxsZbrAS+9KTdD0GJQHE1oJD
hsLhi1rR68qT7johKBsMKx5IqlcJa/iOXUwxU1nsOGRQeXgv397GzkKCj2XipfEg
k7ceqDWSdyEskXcOvEUZdVNXfKeNBo3Hb3MXvZRavDAc/z3AfKCPGahw1k5IwRCz
cJX354rMI8AkI+azO0r7MIQMW6uRYF00t4S5YDFDCdfcGsJq1xj6zZtSaB2KMtJS
fGB/KNVyExAuvYpSi1rSXEt0UZuM/V7y1qJNr6sFODT/NcKMbR4/jOW6ZqECVWDM
A/m2j1GKDpJTiotxY06xq+pArcWPagwGw7RmYYd6RirjF9v87Ih7mPt5ijiQNKCa
wcM8B7ZkquGwqJ4qbBCXMpUIlCSn2LxhSq+xMolIMssYFrHsK+it8Ywpw1coML6O
Yymx0kTQB/G1t5nlLkzIaTtfLNJqQQC7G+24diJdYv7aY9jle5TkvHRhYsPlZj+u
gJKiNX4Yl2jOY3q8iEnbV6h7O5FgsGbZHn/ZScfXpzJYCPbIw0jfwaj75plxy7tS
BdUY6bE4//tI/SsP3VXfVfXy+sVuaGFwv+hhvKXm+Cx6YC+8Q5YRJ7mILrrvJihi
3QedmefrSZZMvjKne3tTBqj/u4Qt+ipiECEP9W7PbcQb8sQISfpnb6DD2hagITzm
kZFKKC8q5t/mgfCeu2nIEfMLZmE+lQs/oJW130XtlnTb6mD0RDaTIRrz5Jv/iKps
BvjxFyRMCK+gaFDzCrrbLTvrcZMEz5qzrzDWXZlsgYF6m5Bd89ZdayVz/9YCftBP
qeIQhJFyQAYTAS6Q9Q/RRgasApLr7UlJbnRZ8mrr3PKMKRNZOVLHGg7pVwq8hKjT
rmpN6rveVlAjXLxgdG4CiRgA0p4pZ5pxF2SctO7Z2gxr68Xv+qP4+guGam9u+2Fl
0OMunv0WM+VE0gtIg6Sfz80vUJFTdi4Rs6SZNisvix6Y5Qkzj6zBpONS2AWzyWGy
Slkfk2AbT9j1XD7Lvk4ZvaJ0tf2BvLWCZ0OnDZSdMTeoMuIpaCja/7fOTcWv18OY
7AsBFDPff2ooXE0VtTqaxGieAybK4ZCg4fvhLrc9mNXQ645L/GslpFRsHSttaHyc
29SR/6CyjmdnT6Lgy3dF6FjwrUYoUykEb/UDw+mAw/TnTssNUbaJ6KFj2+kjvOXX
cu296T+DuvMCEwMFa4j08SZ1PxdDh4RNcGwkxDMdRH8R5MLp9mUr0Q536AY3fr4k
7mEwB7bl9Nw41rpw8m5ARf/Plhdjv7EjTAFHavmQ9BsVpNdRnmd4SkHe7alm4Bd/
Jb7/XX+YYupLfo29P/RRMbUDdOTJu1mXE1ByhTk55aGmIwRiDOPNR/VSVUNho2Zi
8sUqHqNdQtwxjKpwO3sIYOSdMKnE7UoCHprK0RK+lfFoQw5CKm8FINfOjlsasMrV
YKSxr97jNk15B75uRRI4YMrbOIxdItC8sA9bc4sD8RJt9DVEyXxJypjIENJxinnS
uJKL6DSw8bYHdosyUOT6I0HJhalbOCloJyNMoJdRcMBKqsX2LQ4r5i2wSrPQgNT2
T5Nec9S547cKHuqBKP2Y+H8JFDRXkCiqgzckPcxzdJw2qXf2ae8QilF2Sul+dR0r
AnNUlsAOwKTuKNReytGGWUtYowxBT6zCaRFp6w/rFnSX5kLtBd/EUEbbGKXx1x8V
cIaY1DdTnhttRCK2OOIu7kmeZ/A1sePent4QmsVXdEarZZzEVt1KzNmErg0oYxCa
ioBUzXRj0dDWP8zi5tDICopbwu30HocxSzx1lSNEEyxGc/2mCDkrstQKZeurgiRu
0ohR4ySYXkIBdDbh8YMA0RU5xJvPZ+p8Gj1LvDy20pMcgW2mFA0bnDdyuzVWzwRr
nQCEVxUAtQ2yaxf7EtEHVSOztAnXZzkzGDgXPIIkaWJ1TVvlY57OIf5QIh0qY7rd
Mdfm5wxdoEVxuoKgGplkcVGa6hvZonOwzxGgrvL7ZRRptySbT0wZ0J56+noai5a7
WBZOquBzyG3A11OB/KykiGTnnW/aCb+fZMJNiA0x9NBDLuTMZc/HYO0nqYg1lTCC
RUeLp2GAOgHKa5SYzxZAXUaCq0SqsfYP2bsLVdZP+9IkG0ZUB1BGkDJ25PFuXIaS
hwcdrm1s0bnO5I1hslKs9JGypgkqUTSlbrjKzV/0OVbHvtNRkWqG2n3C7TTuuYq8
f2lL3UsRI+Vie5gzhX144344cEgBMfKulH/I0ERRh5dOztOvsofDtNAhqykg3icq
2tM+MpUVmH7n7ch25Q2RDEtQrKNPmT7cdT742YsGpvm2KqL0hZu/K3CVBfVKHKdx
CJVS+mOMpryNsu31tZpGfxrQNWYisi1opMMea1oJwz8XMvaXZo1Nr1hVjmw8mBD5
+cU8ZcBeMgYJVsPSuSpOuYOjwAafazgp+55QX4UUzE8AOLgK/LBcouqiLDr8Gkdo
dXESCgES+yoQikJLbobibkQOpFE0bL9/MvORlsJ7R9scx4wAG1k8rONChSkmONt9
qJURBHFzyJFqeOZ/YKk5fctEfTid8uuQQ6qZ6zJKu6h1nfb6Dp7bVIvsgei9qsf7
FBkeXP/HaXzMD7wBGsZKdFwXnp9MLljeRx4wJnTswX/qvwY0dpvM2HxrNcv/thBa
FZMOHNRYPZISytK7C6xRBzxVcyR+qbTlh72noQgnyxuqQuaou1O+ctd35wdUdFGq
SZ5tevY2Vwoo463dAMsBLIunUnPSZvpLhxamQPclnOuGL8vsYEufHGSNWO1fGcAN
qf41eGbZ8FLf6xpTmVZrsgZ24nFv7Ph52p7K5WAdP2rgKNBxIsuic0uijNiz8IW/
sXD13ptHbDADm4LsBVowlI6yZMP2msDpF+o+qzf+sImdAyzmbmr2+D8kBpYYTwQC
AqTg2YbIQ84/S6is5CibcGAbYNFU2N5m1rZsADNrVIJqucP8okF2xgsdhFe0P4bV
mywGA93sLjttIa3xASY83mR2TFBLR5f5OadbR7fwQiuyGzHuEcf4J+aUGxfcNaO7
JuHBHSBXXkpaUWJmYBpR/UxEQrzbHTLuYyb48wXQ8P7LSs6TAwmd6lsfMD/ET2pl
svjgQ0gc5obREC/OwEbFOY1pO8TPRzwgumS5Bz0yrqoSdl/qzvnjnRuMKW6szjF4
po3QFuHzqjjs+HdI1N7UrLdPNiDodxP2Zli8cvX7iI6F48a3H07Eo67qmmkBOS5b
PKsXns7Q3ECQZSfkEbawJZUKLyvwFxW7zqOfK9Gqp6y6/ypo++OOn5b0b+dzEgii
ZLONlM3jFoKd34+E1N+uyhP0V5JPI+X3Fo25Rd4Q+GgXCzUprkkP5xsnahvQ20HT
dSAox73du0VztoefrFh5OpD7luxJgFAYdmuMMF89CI088vfMjnciwmou5+gZ8Hdj
31Ivdq0eaOzWgzIsEDIia81VbqwoAQd6ouBQNNP1DTnOUpuhrfYWd+We5hTIow2O
WA53KoM00o624Z2PKx/060Ft618OtR8/ErhUiaf8Kj8O9bl6MYuRXDEfOJXi6fEV
PI/3ilKmpwi/+7n2A7o3VPceMzQnkex2gH5FspwjMKedH+aS96qyw6vzdROrpf0Y
nCzIljh+BdiQ48CxF5G+DY3Y0k0ewnZWQOzVq4hZM0ABX7WFm9IokkPAD+JhO5uH
Z03ID88ch+huJ942x6t5ePj8CuDmYfnT4rUpggFjeXLVomnKCQDbRvUiYClg03SR
6v1hCapM/3AChttdYuSHZ6TlP/sxTfG20MyWRIDNhVITpgBQ38Ywcg3J/6W41ot+
69UNdWxKY8kBKWT2mCFzS66GZs+Fb3UGAPhBRK2vKwwpDckDMmdcBznfTbXMQtZm
HN2xu9HEIQxfaISGmhtSa/ZhhCa5eJW5p6OWphaIf3uj2vnYt3b4dOmPFvCSY2xe
6SXXHMMsUN8QDVBWQHnZ26t2OacNmfPpv3onyqn1SiB0e6f1OHV+XFylCeCmCArn
FUn3x0I3D+n01Gg5oZnLzgovh2i1ydiUzZmIOs9MpjUrU/5t6Kf+JnkAkaDluGpR
672F0H/pqzF7Lg0U8lYZ7txXtXABXsONn2+yCFL0bWHZGEUb3dhnheasElSq3LxT
15TgGd5ZqFUEgzV6rjm0WzGEQdKMVdTTdTSiS1nUxoJR8FoOnRCDuhy3c9b2y+1n
ysLDXOcHyC9RSpr4ftKNwlYX9H5ol+60d5zV7kTXN0g+vKm6Da0roaFZGCozmZIe
50PCFAx2W+OE7of5ie9M9bj9n22dkhhfZUTTmrGwpEj97wMg5cgP9L5H6LHbZR5Z
Csb8uNLl3B4PahIvjU0w1pRExwfk1Xw59d8M1jbLxyb0PnYQIZR4KDJiy+dE9cMP
5Sowc4KUKj/waZXVClPDlIRA7OBmHwLwuOQm6MgHrgAI1yP0Tr4TiYZVSWgfBsY2
mVaLkSfEISErNSvtwwOm3gJx1+aIicyr8MFG9JawabwWpCdQqwEwFpePO8e1T/vr
HbW3hy1QsFhVFdlsh4qtxULzX1MgAAa2UZ6TNtJa+eCboQFJTwV6kKMgQKm/lwWi
Lvn0loKAZwtTtE/S8F5+AxGBMsIS09PgdpJpwsn1La1L7A2tj7ncYe4EptJDZIb3
uDl/gzSEOGG4D+/ZoeNvZhE4dtzKQICX3LWbvoFUt7IVX4PyR2xptel7e9hNXmGd
kfsWw3t8MTjBEufdIhtuABe2iKBs/ltkQU17wrtg6Q3Jlxc37+d8Lh+9srxnxY7H
1S7GoNHgzSoZe5vGSxdoTejkWD/6bLhu3mJ3zvIiFPxOcoCdD07oBzKFoliOx6G2
SGnhG5sUetMYwgYZ1qBjLDusRSTbSI9dgRm+cMzIOTBQflAMJ1gX2rd760ERDzo+
RbhKVC7ZgIh4GyUZWQHWiNqg6FkTyYqUG/uvsVpacKdUC/htB87fPoOgnW44WziR
wZHEr5W6lQpsIfoqRkq5+IUC6wd0YH5mctbYWIQ1/LA/x0PyeC7iI46nlWmgV9pB
p2Ie9FLXvuCaXvKj3m9ijgWgZJUEhjZI7+ELrg+N4F3sGFu/dSSXBF6QODoesGPi
KXlEllIHVqAvs7096yiDYR+L5Ah8hSq6CeiZPjiOWNLYrM+wWPfQWYkr6r4vlK/Q
CQJKMtObJwx5JsL8XQxlZy3398PdnJBTv2yl5o0bhiu359A8VButDeTEmimZCU4V
Rh5tbrMTfuh6CVv/BI2//kBOIgITqt2AhBCUGS3zgVoGDXEgVLr00StlMD6RHHW7
MzjwpOmWlWS5HJRG5dMzxKPTj/Vq4OclC0NNi+vCkdgz7EsayLCoFPPQhCdqYybc
CUXtdVqSANd69gP3rHBJPi/tz7aC/AUsHIJe92GT4rk+yJ5W8nyzMeCoaS90Zc2e
5Ozz5cgy5k4+DU/o53K9ysIPFqqGhNYl0bIp3iFZWcEgJCJVQ6r9PyT/EMf8Bmgx
w9R1CQs3JRA9b4tjAG0PhX/YfyarqCjOxeH52d1d6xE12Hvn/flb3dNcC4GQKdvC
fcKcbjcv9TK09xu/H+anYuRJAorLM2QDb5OrMzP3sCF6vebGn3h5agL0AoPgnAt2
OnUNEALS3qRyZd6NgrhhX4tbyXywzlXbuV/IKw1pJCrY6LZSrI+yVKP4N5v4cPUL
tYnwbJtUsLlbmAMgCBlQqMn8oTznAfJcPMRhsnKpYI52qda7GNnpAprL/LpRFKDj
YRjt01wYvJA+9dPb7DyEo4STo3L6RVwzkVm2IB/czsrwLjH6TlPMwk3zXfKjkTLB
eQY7xOksGt60F1AKMdzP1seV8ARt+nFyOP7MWzzFVuyez27TtiBShoUMIlerMVTo
gKJF6F6jI//CzuNq4a8YKPaeHzq9V6aC2WgRVwzT1ZfPC0wWSBX4alYtFWW+AKjm
rmEOdck0/l4GLPIZuG7o//ud4DbcI7gPuSp2wP7lNe/T0wpF8vwvvOAm5mdG48CJ
uCUXbo9FUyJAa/EdGFSmffPb4iQYhePGyEpDIliVJ436tmFjnGQLS15Kbh5U8RuR
8jrhfxXkVEi2Q24oX0n6e+o9hDQHn7kpznHdW65wKmMMok7NewuQqsasCLWLC1GP
ibL2hclgangSP8K3wT8hqq4NibGwuJYbKIEpjuF154tVdIx185mODrZ8jA8vdSK4
RYCidZ88YRfS3kW17LU8vHdOgfyLfTqmSdBL2+6bVQJb2DHMIoIZvezZUKAzsndj
VCsYkLsIU5zmGKYTUtMlrK939adZlRdlYTJx4Y5fakzmN04XHp7mmqdA/bj9svxN
0+0cTEb559l4/eWZPxl02hYTBXdbnzMPhzWnVGmltpftu/ExcmIBzndGVNc1DEKX
ARfdYQXmCq9cHPp7/IkxkRwiONwk9ldTCpHLnW5t8Pk9HCh8++iYyHdexrn6FdcB
+7+k0olY0Fl9ImXCPfCGpFwhrVnRGI2FcNZs5LeR0R7VzQHb5yjeMEdp4uBnzB9R
ARNjpjLcoVZnMsr45oed/RGhbWOD29NTCKWEgmdHtMudMe7sstRduR9/p9LA57Fn
bdCMiASpP/2pnWXZ58PAFhHcOQocGMxossmce6BWpnLdw+WkvZW/4HcS7fKDEYfm
Fkxh2bwRgLVxVHTwXCkAe6lnwkw0BHbUVevEA40ArPigoowl6cd3TlTvSVHodNQ6
6ziMpBY5AoM03+MuajIpnbCgJNSZipYRVsqtjrlA1vWelA21LQfGS6a3TRIxocNO
eYaByCK9Q3vpDU6IHzNgB/Thr7wVkhIgnxxY8CN1YNfBmNxZBgnWY5qXy5x4troA
oNtoZCe1kJy6QKPA+fOK+JyiiHVQtw3f/zain+CxbX0CtkB34U4Dlsl9Oqv2kFTx
phhWLaTBsLxM+MnJ96Kp05Sux9lBbMxhx80h43CMRJfq83URA8arykgxaPFWvUPG
WgUVQYtBlFLA6V9pE/hcpEFfjY4SnADBwPO8l60saJtfF2oyPkR4s6K07/vnaS+0
vXw46lTOkKQL6gw14mVUjSfbLK43Cq8dZIB8ZRTJAbCd0/f/UGhKeLv8QqJLXm5q
QhGd7nYld3hWlovv8hhgbM1o98eN72zQAeOVkepB/gzfY0pd99g/KJ9IDea6uSNU
EHpsOqBZB/QqojOQDSwAEVL1futtOu4Kct6c6enXR5/Byc5a7yveoQRzdCIgryeQ
lcKwIC4ZnEwI4tptFjdrJd6jpVcjo+cWp7IHY07VcB3DSEHX0xnR9rjhosQpD5aY
YiXhMELMVzxKfVqxbipHWMrFAUbazs/DS0F+UjDa2PZjxadg/xEhhKD7SXWwdUmy
hmsj0QPORKpSV1r3zYm2Qxa+pOtNZi/G8iZMPcHe7+MdL+Fqv+lPnJYSasbkbkac
JK9kecGMNjSp2SA3zjEnAHXYw94UAKWG5GhkJo4wpuc/RBbqLNwW6AGhVbvRMsrx
ZchxiouZeaHVRLJXzVIS0CUFvjLrpvv4rsPN0P1GYGyAC6Ihx+e/+Pm+bYxQ0SS3
LoEZkIl2GRGuTBjMXCP3UG2kyDBw3MeZjNi1TS2SjvPcq8U/55z/TGkuvOx4yQJp
8XpJNfXixL/5RBW8UlAg2lNsmXiqgYzLcr5k3ldqeCCQy4A5BukPeDzlyMMiztQ4
3q8MrjJiPFgc+x68FWvmvttpNkTAJO3fqcXx1B5cNfo1eddFRnZ7hXOgZhzI11X0
tWgZcidiZgPWsnWn5YSF+iEDksoitReEJUrLQLCOIujGNDTgD9uQh9bB3J3roQ2y
MN+hvJqGOUO3Q9aCkieZrGb9b/WfkyntOAf1AweoqUKf8Cp3vtgTkmlLelWyU+AB
bDgM5uIalL7gzTgjqPKh/VaMJgqDqz/cFCaplYOAJXEnXAxHHCjW0C4ldZ4hfRoN
Xs8osfdycLQcIMiu/Av8T4lR0f5HBkqrLC988Tl4zFxWGljqx5ZT0zfDi6WQUiPi
fHzd7B+9N77EjLPRoYb/RaB5E8/CBF9qC7WkWnN/h5knG9WHAkX6A5UTrTI5Wj9I
mONT2R9/pDwQFvAKhr6fsffcGF77cCFY67gsKcLKk4QIwBeQb08hp0jAaOQdiUlE
6eO17N3Bg+GhwjcokQhFkQ1R4tZ74VIPX1Nzb5AmFoFDB8zsFtM5LrGs7zbzNLlI
EbUe2HFknArKiZyi949fJg31k7E2wS/MteFmu/HEV9DjHfM/LOekG/UZk8VPnn8r
oqVtpQz2vcphWBnZ+urDqVkPLOAMgXf9kJPtaws2yN5hq69Ksdm86MOJv8ae5eeX
RNQLY/OOrxR9sM4XEfhb7GXuiVmkTjzJzGyYV8dvVgE2zruLTX0Pa17U66hHG84e
pPYXu8kN3yi+CIwkln9KQuiE57US9LGnmxu2oHvcydB8RQ/wMaipuj5O0tPVqqXm
HUWPyJDp5GZtr1SnJD2Bb9xh54mC9467Ck+SvtIO8UqLreyASgvC16hwHMXVMz5h
tw9LfFdfUutsemWRVgFkVpJcNKJh8+8T1fzM4yokn0LxQnkPKV6Hd5utRo4beg/K
dEPNLv3wXszEY23vw3P6SQ+n30Jm4QuIDdABWqYxWv4MLYzqvvX35oNfPkiZjUIJ
EJwYK5cH7kaUGcmW04PZoan+9axSZyArmGw46sm7t2AFcBH3YJz4NkLVJxBmpPjf
S0Nh5Xb4Q0HrEFHY+LKrO07PGQBM1OGeNrGiMZSeRuPmlwcjDkPkolNdA9gBMvOS
vVXaLm3ZNSa2klwCbis74utDWcMI6GI6FtVDe0L4TozY2je4i+V1ERsmVhHeLo4S
t9xT+jdhSSerRheXEnKCpSwTBu73Zq4Me84ZIV1GCgLmqfjvXaz9BNh++IACoIlQ
zndUnA1vfi/L+HcsOoh9AXeplrv8/8jiP/8LXtFNDq0J+FVFrkRZuATm3DkpaIrC
4IuA5jNLDs9O4W6ydAErkczITTaX6zbeEdqh9w1Wl0cddD0R5FuKIbol3q5uJZDS
SZl1YXBFx7CXUVE56hQXLA2au7GaDma+8yG6rHei1GZmhF6wwevPnP4r4sF0iVry
HpK3d8aM6Y9ufoK+OFueJU6rD34qdWwcb/36DlmUsz4E8hM+yPW4poOdU/XxsVwN
Rf6MfrJdw7coeNDo2KAZzKCk9/oojlPNBX/ADZQUuRS2jcsnt05jUawwwnrElAYe
jWOFYILBULi2G5QVKlymauqqcEPVyPrJqWSLBilmVSgTUM6IpXv49bCsYCYC2FyI
4J5bQ70sypCn+Imjo2INKD6FXNyqfbS5OwCUbqA7d3VOIcL7dEwlwzLBzkb+Lg2O
RMwGA3dvBTJXSht6yG1pDq0M21S6Ss3HRa09cCdHiK9/Q2mbAaBQt/V90Kii5cg6
y1ZIZPBMxBntocDILdHmd8FGrmVPndqIJYmlr19mqselbcLHFMcmvzdpIU69pYOx
4a3DvMqj7IAcujabK1GGNaoW5N+laV9R4Hj7lLSEn7npH86jVlBBpokqCAToxzb0
iBh/GK9bErTXs/6xR5C02FluToTpayFrdrO8gAv8Usyofoc9369CYSfLGCQyJHWq
I/LQwYGTXYIUNnElkR+YPmRrM/ChWAvNaxtDLF7jpciV6rB8myDLpgCVyYgZtigX
6z4582mXjy6F+cVCaE4Qg/bVOCRzuW5/0rgv0sEX6z1Nh52cPVWbmlgqyS2Ky0v5
0Pee3qnHkdPbh10CYEgt9j+Mg4xEY9K0s6ZH/XxxI6Q1TtcufjlTwpU9JUNt7kBu
4CN8s7h0YMkY2zK63ReRFZSJrnzNecq9EIgvmD6fpKRBhLzSzxsEYZ8CAmJiHWkd
+uf9XL+AEi54mYlZ8lzYAS9eNAN3fufteYG1FdNdSb1MHJHMaQvqUq0YOY3OS6fr
IacqtcnQFHCybGuXO+nCCzFdfUb7UgUmZMqddoQ/uMGzGFw4it3mXKZHL1R+Qh3K
QLLYHV6i0f/76VGCduUjhotRfptjiFpMKNV//boiwV9c9Gjh6T689MZL4zVSe5qh
DMsDi+YgYys1/kuL1UH5B8115TwW7t5XqGW4DIFR3OOS2B/CQ1MJq1ZJPuYf5TKw
jc//+XEN7ShEHLEf48SCkhwSzBOXXRFocfH55kXrubt6+kYI/93jBN70Bqojeda/
Mv9gz6Y+UDxWVYraLse5bmJmuV3TlsKu55KWeM37CrZIjHmX83sl1eEvtxo2NhIc
k6Shx6hlsNoXCGhz1/blef04yrRP3MTu4buxDAucLmO+Ye9om9ReioWtrZs/AacV
s4SlVn0IrmoBDykCgXs234l7xv84PKT+oHvHkKmgiz4RoCGFnqed3rvH8YiZv2VS
fQRL9JCwnTXPi97H+e8eHTbBMOgqaLuqRI1SiFllXIaZXUH2gm0aOu8AC0671Ekw
hHDmmnVJI9n3ThsUP3YjcjT6cjtxPdXVRdXRmn0cx5GNQ64OUpje+BlimHC5x3Kc
7n2lLYPzPOVVZLAFK05ZZtcw1xpr82JmgyevfLJzekumjrr0qjgfcglsXaVn+fSq
5upiAeFPH8rfrF1S2BfOvaUL8gy3InXK0HVdn1EEEUmQXUmM0txywBUO5qXCVi4a
Jcb/2E4BIaWgFe7CjqCSale/AcAQKSBZAAkofpgMS1xa5U+bqLdbU35lhDf3f4Fz
cVi5UfUD7RB1lAJXA7tB1veCmd2qEEnwzwGJFXXzT4+GqodSs09vKqWAN1NDeTVW
MHeXZZlHQHESEKv5F6SLr0oj2P2U8bRxAci9P3ivtdBlo/EYVvjfYHKO5/d/t7WK
MqukV2DYLPmkHMknn10e5Ii0VDKMmud7Mm+ISCHi4Lr2JMkI1pPt/FjV1VCY+UGX
T7QWUX4k224AAeUqye06r/1elVNNSr+8bv5mGq8r6ohANfsy+FPC0LBFwzQa+WoB
aGE464MIW7SSWsiVGd7V+859Kx4Wv/9AGmngeLaZ1ZmbQ+jCp0xZDYiyXoBQI3dm
F2K1wGvL/MVKsXgMXX26PPec3xaUfrMKwaTuhRsFV2HVc98g3OaG/qXSU1hUhN0w
zKhax4wUg9XalCB4ygqlAlFPN8yEHkLNltTLMCVPHEKMBM7biNCEWbmbc549tIfM
YiPhF9JENaQBRUjNYbF95POis/qX7ipgCBb0DdJITSGbS63WQxr8QA0hzYuXvBzi
cMJzPLuA6y/5Rz7OUH5BxV3nJPaR30zj5ArIg8pHcXcOYLNJ+jrlldkJxeF5OEqZ
pXyZ3cDTfl1zBvJcisycf8IhNEd3LC1HyP9Tw7AqrPJNpgebkZtZ93tHZN9J/7gq
75RxP/rLSk0ilnj1JaHe1kwK73uqaX9P06tw9cFUiTVUtxrVQzQRNGaXXhh31cF0
0JfIiwII3lJsAsff6qrLIYF1Zc2yayRx8JF5c8WdmY3bRgVhVgRDNLNd5lfoeYvM
g0FMaXyqyq7W8ruZTv8Lws3bTYCl2V3PBeHzsnYm4UxiHMr97Jofs3StiWMwIAVV
krR4xKZKpkVa33VKtQzVW0TcAxEKW2Vsu+OtY7DcXoNBqUjnYjdA5fd+edsHZ/Ls
5nDSJqHMzLa6+Eq6AbDOdc41w25FXyUYmnEnMmbHSEH7WTv/QdFliPXGFKiryyNb
qsS7pdwF46D87fS7zKAbG53IFIP11HSnAV3GoQSqT/+g8ZcvlgFKvSLdb49cw6y8
I5tVejSi2gw3Pd0nAbukQwv3MIXo5AreJPZbikDjlp67h4i2XqZXLQu5usbW3hpm
TgVarl/8a+Si0z0LRcRxeFyIJ4eumZS3QbhRsYuei4A/fluEl2pCINq0UstqsivJ
g9FlWvKdmmZpGJJqa2KI9roti741/Ut2uCLC3VEHbSB+rtOjc1+11SHSACuU0kaK
s+p8tLAwWWcSgIXDXb+2SWHYSwecebaPi3ca8LpkNojFh1zTstjVb+lYIZtXQDAf
zAjoMQwVjG6+WOlbD1oPfZhVqTiE3dTLy6nXPo3XshwUa6w2zaVwWJE4+V9tAADN
yb6ZBfVwGNgOyeDqHudXfN5qMnfN/ipUanevYSGCYX3Q8ZZ10qjTvyj+YX+6cBPy
fjD+fgPz7MduyfgeUYKUACOsEw1AvTJmQpW05p9fyyFhKKonPfn5O2p8/ylN6GT6
uYmOEzt4TMS1afVpCy+ADd0+efD+Gvse1qhy1XhzaJPoGnGIXoXo7mHTUHYL9mLr
/ltsnWw1qfnsVSDxB/LLdBDYqdPK8EKu9P/OsFzcmR5BZA37tLFHCXfYe2+J8Q1u
HBk+XWubFRUm633W6ceV+KBCKjpl8SFYwZNgBar1xrSxgcOw9TbFN+YtMwdESmbU
zsNRw531VGOfZx9IGEAoTtMNh2AVFQeU0Ba6TqNsrC7ZJHzjIUvbYWi8OAInvekR
RaH4pUZjVA/Qy0PA5wUuY4U32HS/JoCIflMl/TBnsou45cuwkNv7XRjGkpTOOmzN
nNKCbeKWlSovqECXLfu433SNn41qOek6t6sVlz6j/RDvJpAJFgn1rA719K4h6m2s
gw4OEiGp09KfperKsu2Beu9GiBbw2GqFYe6xBK0CshmvR8TzV1UV7DlB7x+flAek
O4+Qx8fPDVeSqfTmX4w4sr3RTSfsncLzgnmf/3o0M74uqqWf1qpAkka5Yc1cOEeb
QLh+Fnf5aRn/K3go/AAbQ+f+GPZhCpKW/vCVN286ISdJuoTL454melgoYVVKXFnE
AngQcYOa10z3DCBHTuPmmq7EyL9rY8sD7vlqNj7KA4cmqbg0VBeYpMtjainLG2SP
VZH21Mu8hPL1mHhVsJZJ5gBPSOi24Idkepugxw0PcSE0cDkh38d0l//mxIkJgCxi
lQ9n+w2I/QzFbpJ3HH7PrbMh2jwPh+jeMGbIO3O5V5kzQsybcduO19mqxe+O6VsN
`pragma protect end_protected
