// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:58 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zy+w9hWvpEFnXHQ+G6HLrztTnJgvhwXG1QxPg618800dl6a9NLPECWRvwCwZp203
l6kjVHBm+ITRaq8oHu5XLoT8jaIWT5UlN47W+1vCWgWnkt30KKb9AwU2uPyQJfCu
+AQCcmApIxiaWvV5LFMhsA0o95TgmPmcwcqqFqnridY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6544)
I/wvcZjXSsldBG4dUvT+R7ZZDcoilhy59vfY5bptxaTxHOcRnXFsUNxYmJVO7sJt
vQGWZrSg3LSI6aOPMGlqfbVfU9SEEKOg3CcizgEGkr8QW6WPTq45FsODK507G7Gz
AebL72g8bpEiaZHhkM4/hQet8cExUVswiBWa1vIRiEahcUah0JLnQbL587jcSGMF
QtaSMx+mxefhpCS0KIJqoOOdwk4QEcrrs9nTZNrNhsJbnmIPqx+6EJxzc8k+YPzg
3g4+bDmzusGAxfB0q3VevMfPwQ5gdWJrWfeFXAFk42HZL5tapUzQwIirzf8O72YV
f1T1C1duRSDUFkH86rehYXitvjYdrSYAVUML58wEo0nKCk6CnZgGihpJ1i1m1Dr5
F0itNAoxCD11kJ23saXLQQaGb/6FQylZIEmLzjN0meWj91LA5kTVB4YCuYtwuBu7
nF4V++Qt4XAYc4oPHBCTmaHSYIbSfn0D2Tif6qUgNE+CPOxohsDK926oMXtenGm9
8PQQhHXsq5AE52juMhqahR8uGe/ZAZWzGLV9jMJDDZANvh1LaErLOawlx4IRVkWy
Zscgxa+SS0jPMI7qP99+NVgBmsZCGzsqrbXGHiCKVrHjmL+2fUFnJV8tqm32zl6p
Dh2vH6yS4r8emX/hMxbpjNd33ZoATtv1FMDfr9wwYTb7l0DO+IVZwmd68ss0RUHt
Oj1eMSOipeOQkzRWUeAIgL6+ltngCbMs9caj4zJdkXrksvaMcan/XLtXQIPwgq++
W2VEPvBHy9hu7c++IBYnvuXIc0Tz/R4efirZo4QJN3oC0a3OesX376COSLsLoju6
oxqIXkzEjq5WtptaiEPqPaqYhwwh/7YTeRkNq+R2WUiV2cYE4+uUvhtFpTvBEGwP
Em2tZoA3T4is1IK+MgVc+ZrjIgcd+QGRy8OnN2OLR2DgULt7oUgvTAfmseI96FH5
6Daklw4eATVm92kr7+4WB7t+E+QsJOf2yB0RG7eXrf23alC+H77TlZ3TLfoaiit/
SO28ne8puo1E6wumikkIsAtUlX2mTvZzP36YdTimgfHmpy51eLvl9d8ahGWti4Vd
DhFusoKTqr4UZOgZe9JlMwCoy0W6ZuRIxwvUea5DppWrmAc9mm1EZnb2WV9I/ws7
CszQg1f5Z5g2gkGXZ5akhoTsHCjtsEvT8QzzxAxhXkylL5dqJJL2f7gTAEU2j07S
Kbz28xqaWK8eIrYiBnjzOuBoPYVKGavxrGaa+BJU/paIIFPgSrUS7heHIMQbs+Ey
ojB1lq3pSCapxPb4YLi9Hc0wyo8MXI8r7hOzUme8HOBBxCxo+4w8eIMfY3UEnYFn
3EEOfbXo7UD1AFuntyzfjqB54oJ8Hqm0lCUvH6ni+rVLeEeHJSoAR2qTd/6OYOg7
SfrVqT+wfNcp2lKEFyRfHQnuUW2gUDyF32j+fuUchnBpkEEq/xOwOuh6GqVpDZHf
qyhtWJ5sYNAVWbij0Cw3YKjVZiInW1u3H/oQSIASOkEOKq2N+dywAhqnVl/CpFUE
zASz3ruvNqVIj4qpiMY2NAmu6q3d2WVCN/4nesI+awN+tLhzVdRNHEbrOq5Rv9Ne
TLUg28kuIenzaBQVpgMe6w0LAJj3OrWmj3JYtK7S3xioydcIE1PZC0wP2kM2u4WH
roLC5GGTFvQ4Ecd5EryMarp0imiSKkATLDUuERJfGjoANN3165Wo5lB4/9ji1MO0
+Kdd8w6mHdcMA2dHZQ/kJHJQNCdspyy+FeVB73BTnJH+oZVuv/43Mx1+RRBcT4XS
/Bp273F3IXT/CgM8Art+GHuK4BA7PwMrqwuw0zGMXy8yGy4fEt42V12SodmztP6z
VP8o8XFgACxNQlaBw9F7zbOmjlP+rnvcSrrTn1WMUMbGCHtrgkdv3AJLqLfqVKvi
Z3nwgO4jwLkgK6yOnq6mcYgoA/Dq+Td6imDY8AzRcY30d47toNOevmBMA2lJoLSG
U/14GhOyl57xFbpYIxyVrhVqKNyKhF0zIE1PsgFKcA2ZJKyZVSGRt/VLQJ6lLquL
Mdqmm943Vx+3j34ZaWN+/Ys16kWDY9YL2asSBi8AokvW5t3EwenKYr8hF9euGW7O
NbmGLrAV63S7a0t73cVcR8X7xDyRqYU64Xc6TJPhozKIqxsesd3JyV4lTcJ8cVy0
TOx+VpEqYAhspO7iaSFO4TrYpfhZty0va7GxQ27sw+f1mCbFp42bIYjOw/+u/2dh
R3e8pLbNmTLZ6BiBBWxQPtzhy54AGZdnujtvKqH6v00Xb7ZXE3CZ0qQHx+RRUlDb
pLHw61a4n6MmUGxULF+J//Ti52TtyilMBHm8BOYcIkyz/Jrmx9tXkjY4JkwifwT6
B44Qi2oYXHtUsp+3ilJUm/dcPxWm+q+8AzNd8tJ668tK/Ny0l4t7G2mI+SDkr4op
ggFtOzS36WA29WDyAm+7vVmUbO62vrBBpZ4X8rVj69BVip2VqY1F2S8yvuqGMDhw
qxCz/tsXDsw+1tHDKvJ6b9ikmyoRG337Mxgts0qtYbeDIYXeeFSxqM6ZiGumwxrW
z87pmuIZZLItFl9kGM8phPaJ+SobmKzw0q+Yt+FqpIoiReEB9IMXFNSh6qYb5C14
P1PmAPFnhqWqBDUzshcjNr/WRt4hT9l22sGfUt8HqRM7pchKIuWtAIV4XZ2msQzZ
Cvbk2tFIEPaRiVxVwE/qofbgWKxthM0/Ai9IvAt//9SgRO+jygFtOWeYyNipGTFx
1VW6eAUOfiVfKYIiAOMhk/jWKNReC9/uewzxdGPV/qe0svsYw1bsv+i6TbTgOE/k
9pfLkRfvGI+76NSUpc857ntO0tRSxTTlIg4fKttCA/I+xri916mdsEVLeG+YJAOC
WZM33mV5JLiCyT6kdFF6meveVUo7nGu75UQ4htuBVduqevsUHVGSQPp5E6Kiq4AK
XH4cGmILuBr4ZLww28mFP6eHhzyMdfAinh5KtefGd98hwlGEEB2sFSmDwz/iYBAi
Ryd2kB0hpU3JHpzfse66AabjWqKToCmLDyyV4sTO0q9jNGs014gUar9BYgejC1yY
4eQj1jDX84onhnmsvp3BQf7wMtLq1d2zBNi0KtObpJLfOV4xp4wpsg3OgqV1LHl1
BoigkSPlnskWMVuvW2my/h3X/wUlqw2PEFgvOU9I1gMi1WR+8m8Qh3I6DwQAfI2o
7zJYxZXYPnVnNNrrhw11yOr0jcDOo2WtBQfpLJGvRmfsbuZbn0iYXr/gJbRnV8wG
bgwuMHw/FKebi8fvOeS2mThiZlyBC7OBoFhqXXelbc2rZa3FB91lVYCSxUJsYB59
z0h0VvAqb655q45IFyd3QJ+2I8CUgJeUj9Kmz/9xoxivDuHyVstfb+VWEzdGXBVJ
c/TII7XWslgVD8CcI4iLy4xUGOlgRHLcbhra+LJ4GLqdn1s8vDdeB79UwCSVfFtg
8ucmRZ7Z4qZogdxREV2Y9pozXdCNweHN5KM4UHCNvBjqAjrwJMPsN38zZYdVXqDI
8G2vszlRyeRnu4i+DRRWq/UfUTIHdcAEmm+gyh3gTEFGBYu9WS762oQnDX5YU55w
lOkYd0R3oDKpnCC4gnrWhFUfFEUOpbaeDeXGeUBT1EV6YKc5O2JId0F0pltXSVGj
zf87+RZ2IBTwi+tqZmcbZ2ZUVNiy5SU0DX/jwSvQoXxXLOFRujTW77gdsZx0MxPb
XLW7XDymtQAvMMfog5Ok5PL8R6XwgC6KiTkiydbSTkEdNeW+2DbwFbKI0j1gHwHa
mBIx98uHmjdrY9PP3IBl0Id/wUBzDrTLJKzb+SlKcbEt0F2iOKGzJ0ONuV78cRUc
5mRizw1wb3AEREiA56UKHDsBY5Jtx7sT+oxiWmIABP3oySyLQDg29hxkl6NRmHvw
zQQH7YCj7TpCwE3l+R1uWQGlCPcsRwRbsvda4wmI39RUQg49yrapkErK/47gL2pF
mz136HHw5G8DynzZ2nkkVQmcdm9h47bX6aylxaUFkhS4xmxgsVHrXgRZu48O492R
6DeH8vGxBFyT/LbwhDYwv7Re2N7vSodjYo6c/Mgg3mV9ip98CvDutJssegx2afSP
H8CMIuZVPd8Iy8Ll9sWX1S05BIIxgNMq8K+OJbp2CaK+dm5wH8vP9Wzm79P72DOd
RGl/7Dxlc1jRDtQlRiK3pbFFYYWsyR4UorEIkYBVILU0ONiIPShwAYAGEKdPTI5Y
9nyTRX0/l5uAoIe/DH230rGPv++KwVJpluIfd2FUjnWWeagFMS3rjG2UJZeF6qjH
BuLid/YgQ3QFw0ZJUQER0Q44h0RRIpImW7U2ohDlpI3X1qZUgbdveDILZhE3tm4q
TVygT45Rvp8OmTnCNiRKmKWh/HFpxwtKmWO5sfwZOMOd8R1sfNRPNoP5kKV3CkiG
rcylZxvv6b/ksQerOhWxvqAl28Ptg/qgwcnHN3DpHDbVhgaZ+6GpfLL7QaipZnB8
paCq0KLG53093Dn6HvxjX30OhXI/ZRnl9xDIbXFaMd/JMU6i8tncpHsNsH8PQeZG
OyoI4GnQkhfaRs1fu5LMWJAUgKqRlK/JS3WxsJIllCizLXzcBpiFly0wBQxfxhlE
Jcwdii/dn2rqIUViXmWcy0wJY2VDBbzZi3ysW1kA+WNfdelsyTYGuf/uMkKwgOH4
EDCd7CTbyzhE+wUi+k1EAtZpAOaqjq3BE+vWchb2uJoWDBy7g0bzSt5lxco2JG+h
GJ3GPKaBlZsfmqozE5IG3STF6wLL6VZqBN/nUPP2muC7UAYT2obXyEt7uBrCTx4B
yzphhNjpMNhccHXB4uo1QHBdZT+aMDBDT0SFG+iKAjvIbOg7pj9RfpwJI9NnC0o3
G0yJVY4uERZ+BITzzrS/aZhZohN89GzSNntFhHndsekmAXNq+VeU6bbspu3OIhFS
HOafD39T1Ynlp23tDC1Ltwdnla1ntXnGOekd3kmvES6XNFgaBp0wYa81JrggZGtb
btLL8SIQ4/qHvWr6IV5nVL3G8emShoQIV0XdGhH96yEc8N/9REJM8QlIPU/WHodK
szE+jryvAfHttkZEjR8t41uTzwoOQ7z8YI87H8+a8j07ggn+xbADGrF4N9pIhda4
c5xhHZPswznDjeArCJEGUpCmlbm0ERU5mKqArStlEbswtfj9WXFaT0qDn7LR+VxD
5VZvL9mFfoEmzBI9V8pTcQUWO1L5xZBet4tvZu/s+40kPaoH1co8DswMBoeiq0jH
AobwbsV5F5wHMiT3/uh3CgyIJwBcv5Sqke/mhPgwb7tzs2fuD+gO/29sS7rs5vPM
iz3/d3TWPGz8NyAEwnjtvlG2j4pmnhKIC9W+WPAw6qbHgEVRmgnrhgO4R6WKUkhq
jLSv0+xkRaFRDh6iE0MCelWawS8PGPi9kw/wi40tYfD/hiO1TAioRvXFqOwqrhtR
AwYaN6J0A5XrAXr7xw8MlCdpw/59NR3il8QuMyHla9Htc7bWkaBuPK7OppwzF0ys
Ez91uvpT/mFJzZBgDng57DL4U9rxxAWztQ9UDIRKo/lkxLm/pOHZOKrbDllvrJvh
R/xvjwtHrkYezAkE19SfYVdgE+6d78Op/+k4tdOGPmDVHMmGdu/dMUgzxZUbbf8F
MtfZl4xrHj5gDiA25yBqAzVga6Tw8xgQisKD3A/hstSuEgIawo7s7an2GYC60Ly/
zZAJo/7vxbbXTKfvuEbTU9ezbzlwbhcJm84//0ebanf18rBdGSIwTOAaXpNH885c
Nu2Duu9Rf0eoRh1vDjZjjVUToJ0p2Pg8dt+1DbOhLDfzkOmuJXrENyLmfkOqQRo3
TuK4n+sx5x2rhhMwSprozhV9huEoWJnRq8x3UjZ235kolpwku043DnOG/b5b4yvA
mwm21ulTmSN6XgQm01KnLqAD66hwZZnuNjyuBumHAL50h9aApbdTjHeFxTA0bIv4
ZSPxcPK8vCUMFgLFvjlc8C75eQmNR9oXYCPyJb3MObh0hKqX3sxtR6Xb3I8fiwls
Q3bj7Tzl0dCOqimsAmmHoAzNxbeQIREROHq1RO5Hxit6Pj24Dua53lKGekDoKKTk
kgdn5hHQKoX6vpT/puSlUwpyPqAlk3hkMgiH+cezMg4jrsdxt05ioqo7iT1GCwIR
sC4LcYgjjPX6O6MgofPXxbolIZjYhxsdtnua/Jv2gIZWXu2jyHIFWPFlSxtjCL6c
Eym1hh1yd/sWGT3hdofMZFAIkYxxIuiTWkthR/FQ5Re2fvu3YrY2NIr1Qx21wfte
lYzsEtFroQoOwQYDYHKMYDANXSFVPlLO/SBRnizq/Au5SoIYBG6wLTos8WdX7Z4r
Uxqr1aiGqMXjz2A1N+S0M3KCFd5JVuV6cHq+v75p3UxU0snjJhN9X2NmXRAIavTF
b5Z2XA/ofSx58lksxoNbfFen11KTYKJ16HxW6zZ2DvGMh9srfDznXtoN26gOGdmy
IkZ3o0LhQy6P+UOZ97NESc7jvDcg+nseR/h4YcjppqdcDzAY3Hk/qKLhU10f++xm
kxMmSr9AXQWrVPRpUfTutIeHbiw56obTRRKgfa5aZlnXjAQspGrIf2d9h4QV7I2O
MOn+qfZ4EfM2/XLxrYFlH9ONm8IC30d8kmidTMEP6dJPmUkRHHmEF+wtxLPM7wnR
NFQk4jb/euGCI0X17dXkh+8Yaz9MU+4MoQmmiv13mgZBbPl9CSZ7kXDam0YRzTVn
KOZ1Y+1Q42oCoENUydoM8Os9n+Zw+ulYmdsJxUIIxsT6xJMpUFq8PGapysNIucXK
BIoE6HZ+PohRE08a9nVJTF7ZXTRsK6FP94jdEglZgr1lWhJ9ufS9gLTXqxI8NdRX
Dxd1FInaHr7P1xDs6m5sJ0rBH9b3/9GQOoLSPKpttzZi31AFd5eCu4tzEMx7v9tn
JL8D/rAQbxeQllXovwBAMGG6CixFH40GKrjJWVrDyH4qtR6ZfkFTSjk1E4wwd+fA
rryxvYXmdTfuS0YNEevmSE/o2RkWYqknev96INPrvMkQjGL0PcBsREZF+BVvs10w
7TLBnKyv+x5zgcT+T00zfe/V1372Vb1bZFbg8+CczZQcBsMIikg1BBgghpVMl+18
HdBQ0xNwmyQiMlJVJ86v/X8N2IgEGuJsI8twt5dNMD0PgS9cX7JR16upQY4I9BI5
6naM+aGXw935hxfySvW16RIewDdq5fk738CAY6cHPeI+m5VkoR8z6S6QMYbbkjAc
mEk2RQ/5zLUYl2XZxgfeBbDOt2kFemDHsXAyYPOak+H5D6r4fdsLZz4Cj8cJYAyo
+JKbEuEjGHrBmyHhsIjPT+/y5bFiWKkTQ8LMH9nM2McpCRAAXKdFFPOYJRzne/5P
nvv50Yim9Iw79uAcKDZmgF2BUsMakPuRYdDzrtDSUFc84y5R5HaQsluFT5K2g9Ob
jEKjSWzNcI1IgOIira1HaAjqhMboIuPKlDrtGDhp+KRKK99Ne2YSpf4RzCPAimXj
6ew/TotU7F09WSnRemIKREdB1gWR34WxehSeuYjjtKK1yiu4uTtcxwBoJzwmBPa4
Iln7QTHB4ZV/GFdS9bfwfbF13qghx0TrnNiAAdRT0XoU4skfP4xwdbqM2TdvaByP
bvwmXZ6MV08tnSn/+r0dke/85Ob1MWfxjLBLM4slP5p4xzKundwH8n7365O36hDv
5ZfpFh/ZKoApiVaZ9ZNb0qsJ1yDZeVfJdF9qdTMkp/33pDMOlvYpQcmdPGNXAdOl
VDM5hvPMM14a8vUJ7jbIe5tWecoleRuMJuEkiV226dJpgbrbqtVXZFnBcxxxh9pS
TPHkczJcEAVkxwcvLVd3gJCv9McLvrFVn52+MDSohvki7cGA/M+uqLjjYJc+tjGq
3m7fOpWWowpDzgKK2LX2WC4wlyZGAIIu/Dz9ndTPozuKied4wD0Iw00BvojxI4/k
hRydTLNWEzEXvjVAl11rJUg++0vXg2Vdcfi1CdHMdregXiqu2uzQrqDxzn6TViBD
+N4xWg20fFuUgruBYG9uEqbCy0nCpvUBy72J1N14T40iMAV2OEDzQCdQBnaSMMwI
TslAJmiAIJaidATIPPeyzJ6e2AADbGMxV+u696jpxFmsgLli8m1jRccK4Aeg2u7s
+nF/IR1AIreSMvtSQ4gjRmZmCw2D8Z2PDRXs62Q8E3pvU24t0PphM4Wx9mGFf/ee
LiFcleTrkvZPNDmStp75iz14lNc0iqXWVEMBAbiGhQHCOMO9d0iYvKvxVRX98PUo
Q1p2z0kovQhnzbi6A547d6Lfo1jBsTWcfSYA7dlalXXWLid4osJoA+ekcIa7WUVI
l0j4p/X3HQ9yzYgvXmxycNxCZRMheJ3X+A05ANr1gfOjGJI6stGKzZbGeD/ulk6/
cnbgcFT86jz/j/cyaXOxmhcaPsTeBywbPS87FbCGIrad7+5SVhzs5ipUNTqG2GoL
JgK3+2u28DCwVU37WiYfA6lUJzrPAozSjT3VJpUZVQl2dhdGXMTWtmHSiezjGUsJ
6JSmO77qtDIVVTFMUQG2sFJ4gnE5LI7a9koJmP7VAx1BzJ1wzJknSyeBlfH04bnQ
589jvj95k2e/Lu40bRqNnoIrW414shYw76DBnOdhUu5cwUXymbfdw6HUFM8HUR//
KI9pQIpuTqDUMNIAyu3Qdl/npPMlCVrEPSQkIJoln5CgF7jI1ZUNrKMWuFxtCfdg
fwOnkr95wO6IHeijzMLEcA==
`pragma protect end_protected
