// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:43 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OaqaHv4JPQk88hpO6AhPqvc/rmP1ScA4NhHaa0uWD8JXM8PTvRsZAPaojqoGtW44
hVsvDHvMvfI8q7ZUVVsjz6aSI707BzOXeCUvmelLiF/06IYa/cEapDd3fhzwWcKg
CqSQ0m360LthHznlE0Dgez0usfHPXFP18bMA7G76vFY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5280)
XTHCcQhZ2Fgnhxw2dQnmLjQJLvruUjKog/9ZuI2aWflP8bmmwOM1pzlzYUIleR3a
NNpQiZgk20ya0sdXtiVoeUVrJRZCww2q332LHfjnZSRHV9qFl1jzGR/lPXCzHXa9
9YqH9QmezsCttT1bYWnX6+P0lrjJZknCDVrB5jWqVsKfDjiqtnOsOteRtHCRO4hV
j0tYox7jgt/8p2dIAbaW4MBApHWO16PyoqtwVYnSH0lzyZKPVdRdEJ4tE167nR+8
D7mSTz0ltRQQiQKph8ALhAJFr9WQqXQR/OtXfjp3vvadj/Bn83/O5cE1uZA6lVlG
k28zxAU6vdhIIBBpklQinStADSZSgoYM1gdULAjEpEHrn56OXVYYuflOGb46UbNj
DutLIJiB0kPRA60ugquxTaReKgkbN/4kYtIRl3vgjOPE5cJL5UQzHldQ/l1ehGI+
5XDVOO65+f+XRqgag0uUuECZFmGQ8WPOFU0FpnUU2e+ua95/qSSnvNTrRwGJQhyq
cbld4MshplCmPuDM0a9p9zAdXTZkH7DKFRsR5pq6Q98KR722MxRVuFA3B37ysu6U
zVT8y3kYtLQjO1Vo4IyQjKUVFbhuNB0z6c1UR7v0ka3DkzjuDajO3aOkSfGrUV87
7uuge+5HBa1jclSlZqrDlywpZf1SK/49HkuNJHxTHWVIHZaYmAemCg6bXqKy498K
DkMLW3di3DIaIutk0BudKVm20cUYVP0ISTbt726vhDvrJljVt9MX7NYvahJdsYlR
pOOPN+3Zp2utC4eBM6zwmoU1NDVx9uX/sdd2BXmGQhgrIhtUYDG/VEw472OOovEx
zRGU0qUtLzmYh/u0enqPHGWM+ctRMEZ0mof0327wd9xts0XjKLYlDjBO+0KQshnI
oHNjR7iOAMX4pRPLnuVLSgwW4SiAg9vXejrVr2n8cWAexn/P2eK3zVYjrstrCa7D
/UMkQqiewLxhKzUXlnM7OpKbFSn55H9bg5+BEF6sviRJdLP7H/Vqw/vXY778S0gv
p5sSJ71MQhS8NPIKLa5V5glrPbVVaHMIHr3aACcOnwiNmTXnXs0yrD6jNNXRbi7a
MAoqXgBuRZ4pQd50qrf0tEYxsn1NXYTivarOvC6sv7AKD8uAKe4f1xV3rtZvYwKW
pzAU6EfZtLtqXxk6u/rK0SPQnNqFd9XCL9UTyrbpqaBrGsdyGvlOu9GjF0cbjKS3
tMnjQh415mwcXeKgf6pydBtoZH3C4pnaMI5XThiE4ynCmoLh5vNq+FXEGDWY7D4B
e00Nl6POGi3TWgFW9RFjARqDxVQaNRHFOgkJn2dZumBYL/qIu1YHynsDPfC1KvQ9
8FYgfHzMUkxTqMSdUwuAZ0PFbD5yEMrqcEuQ7cKrrKQ+tR9B5eJHLhQoykmH999E
eqCi6wMOnCKpi4CIf7g05Ikmya2ffYIfYhE4Lp2y6eFoWlfGfOPiHqRjSnqUv1sd
QFh7DosAue7foM+j6RvtL5thyyfKfz/7JcTQWp1bDwehIcrJ7jNCrSsQmNfW8jgX
Aea/pJqfKfUi5kcOKTFRCMd+J3RVDETEnO6Sf3TEivhFPF/Lok3+PqqQKj/HE3R6
ilT0tIKSFqoZIn6yp2ltp4pnOxHYAx+pNxvKNcsgI9kEzc2Rj6mFRQgE2gzxSBKM
KiDLN/icZd8uPPG+6JDzL47kvMjMi3RSChAzz9t7GhA+YXOB6AyNriRcdsQM7fV+
9EqAFmrv9A5I05VNmX2zdnews8XzgpMXGzClXPSatuNCMlxdRbJSJhvS3rHsJddd
TzPgOVSpYQ6MEruH4KDi/LM7wkJAKCU2jHBz1gjjNjc8XfZ7CI+J6pHi/5y8QZSW
UH3THAevZe+ver/h+N3he0HhTl5P7C736qd42NW3wi2zl/NT0BI3TNH6J0FHIlXY
AXJr8UjDgsRP0y6sWXrTMmI7YEWyHG/cYsGpY3rNsshE17PG8W7lDKyaDCTGuEpm
qQbcCdC5YggLnrFcwnQzdfOExXkJvX4o4aZiSzh72wHla4T3egv7JYkGIOLq2FPS
ENt5gZKL+gqnEYhQoda6JvNSE5Zkh1Pwy0E8qOwbmaTwqS+HSzYmxi/THGaosrvq
pi8uEPM2ZJ9QXJuDf/G9AlV3iW0QTPVDCDgceo86G2WLEoQti1UZdwVS/yzUh1FL
RmUAgEFk0Nj4A1tYgJje4Guc4RBltpPEfDyQymetn/+4+YjbVZP2hYRAjl79TOsQ
InOv+ktHnKA6ORJuyi5jU4KLuOBXZ+i+cZLOlW3Xl0yOkTuWTb9V1v2eutt93VuA
LfppAbipqJ8G4WmrXZIVImZje3KrmT9UUSgOw+s129iNFzheP3LstLrMWVq35l6E
kaAV0EPOLP0X7/zHwJhmgyjiWAkFyOWox81zZTi5Lr9peSTdK1Eb596vhclmiXcK
ZxITbzuzWVbyNPq57ox0FrtwETUaioxNPdsRFt0oY+1mW2P7JWqpyA019iIttVlG
BKeOtbgDfeuqIvrlmWPCRWpB6q3/7uB2aBm4sMmfK0bpevvlSIlEPK/aEyiLKaAZ
qz3tlLRy2/bdsmSKVIZ4xJGvLjGYOffkURUqA9APptzckG7h5h8bmXr53VfDlF98
OOdE8ShNQMgds/KanzVXhXFLhliMK1XaWoJbh/U1zsE/vN2RF6+G4EHPk12laGWD
O9IRyxhpsnZ4HEg6Zc4Qg33zJxMwZ1/YoCtnpasvEv4VW04966kv2PA2lmlND1wq
sW1VWIC5YXtL5NvIkoEPUyN55I1Xr8/jAZUEaR7VaQF1xQWKzWyzzw89DN+FJK20
cAMa9uYnRyHTEikXr+Pao8kIQIkfowBQOHHUpnwLbW6k4829vAVFGyc+S5gs/cwe
Adr0ufP1ZsBqaTgpjT8QXpscm77auG/k0VA4fBwd2EHMWFrQPvCMMwtlqYSoGCQO
Ara3wXR/awIh4X/P8TVbKSEngr/8ETUyPF9fYCFZ9Tmf12GtNqoLDujGanO/XmMw
V2S+esHdLpbNILaRzH2tFeNQRCQVaCSmXM3z8LwmUferFS9Gu7IXRIGUk8l6jDsm
Ybk95KHb793xr1/cvv4ZWljZLIqBipVWIQvIjNIQDZ9Tq6qPkLppkEa5Uev3LsZd
yFBtvM2t50u/e4OzfcVcghqJeI7JbIJ4BTQvbPA/6OgyKHpAvdrCLGOj5ps1LqrD
aKF1T0zGRaTqv4ZwnnRm4Ffd6xtX5mAZ17mHv1e0/8kpdwO06cNXniUg8RuO5vV1
wBSilX2swxjFOQZY3OTIkS+QQlGyfoelc+7CB4djqvxXiDh+q8md2cbMDap6txdG
GQI2XRWK7bN3rap/Fi92/ZGaWpAnMlxXN/wPkFZwqzUOSD+g8oGA/9mnyh6VCiHB
OcbXW3+gRDRvs22rzMxJgqnVZPmR+vnlaaQ7mBALmZBxJlCMbT9ZYtrDNnJzOcfa
pxbAzHQ4H5QbKfwQDXUy3bRyTWfV6UBiEjAcEkNGDWecj4Pn4pt6+dZt9RHWvLf/
DPPQ1I38fzOI1AxfZv5A38C3oSglsHyG0RqWbypbjM0+v3n1JHF3yRxocJ0896AN
R5+fEbSdrlwFhu/bR9qw67R1OFNiGrULBaIOXGBsJjMeoHJ4OJA9CTqPo6jsgABU
4Ft0p4c/M7nS3BrXH3Q479sl5wCESp9JA0e4EVo132v2lUfa5AgBmDFUuh1YT8c6
ULahs1aQVVrE4WNLB3mdn1NIrcIYYDODuP4H4r3bPTHzxE2zGSS/dX5LzDm443La
6BrGDsSzmnjOeLcBuyDt6B5L4V8SKC1QN+7ebLvqqsxKyZxhQSCGjPmA3ZxA5XiD
z6mBUkxt8Snh4ODo9ZKmVsUiNv8F454e5ZEy7nMhPD3A4N8syZUe3q0d5lX2ZrVd
ENPSs685J3AVA6/IDv0NZBtAMyxfQOvi+d9ll1Qy+KAr8IQu7JeUqckts+FKFnij
G4hu1eARMEEXRkMdyHnBYwpmx2VwygAo/6tfINR4TFHeUVeQw4mU8eYyZhWMh6rD
66t8W23lULALF68v/71475fHA+Xc9yV0V+zzQbHSAMkalAvaDrJfAwQA04trlAHf
L6Slj2Yj5okVN3wAcWuTzc4bFJFpYBAqklTzVNEirI4e55R4R/8blhtDgX1skd9y
MEWosan3ihBsx3zzroPfGlHEaT/lrhjD1WigusvR10tayl4ukBTAk96gjiOygQ8s
27+iifuv/JjS9Dh4eibRK0HENBK7aJdnT4P0em+uCPDCQYT4Rc5t963KUJXPFeZu
46YbiPS4I4CtyDvecQthfsav41dYoZuqD/1dlPBT7YMs1fPzI4Pe4JP4xlKfYPKM
yXMM4kuzJR5k9CtdSbkfVjRiT8lBdeDq48iK4C7LhY0LqZzx736TJfZ2BlHpcZyj
VNPu9phz5HCST22xyIQGeH0snzUmmTNdXWEuK0OS29TTGayeCLeBAGioIgbwM5rf
mbnaDzUP+UGJB7QlMlIwENMOkQaeyvudf8VQpHi1WMc7IZed3GtuZH6l38KqNBhz
B433joM1zhQSCC9UwF6fzcK+OHFUxHQJrFbUdc3aamXUnDYZJlvNTKHSEk6LVf/L
/lSba8c3GPu9osNUjZK3XjDbc3Prxd9YQ1A8g/dDroqxwMHMVuTc43b9MBl8SHfO
bLEkHnBPYm/G08F2KlP/ICZnt5+zEGhK6sgiy0ovRIz2dhqo5ImAGMFOimpN1i54
GL84MII7e15VCUJtP7oWRbIbypYeBNLWaXqT2+F9wV6N1b9UvMtwPAhqw754x1nA
xtDZIWJo/poN621wxB6M65ipva64XsAP/8YKxWYz2tEzCjqig9wDKgs298JfEGXg
K7YOrHanHTwNsTZb70r6Za5upItbXjumehnryfDERGHctQ4Q+YS81SoXwAPEFtQ3
pM/iI3hMRhv23M+aBoBij89A7TmAhn7GY59NXI20uhX5DSg6ci2tLJvRQ7uKaZ9I
UJyDU/IzXbs5lmiNR4M5Mz+mWZQjA+S0gb1SB/671JWl9YpM040ehuo7Yi5qZkRq
6qNO650/G7KQLZVUJal87vjNl54R+kZnRR4YVfjcwvfEuLRZvgemsKnwwE3atrD+
BjtXC1mb3yyalHQDy+b8IRgqL4tDLv7L7o4boGQ/SIREQ/gzTxoBAO6wD9aoyMnz
mCCFxWe+0c1RASYchu26vg7kBT1oqnGZa8Z7PmtFpbeVNoglr+eNwrzJW9N0bYoO
01V73F6a8uZbTOi0OnAe9sfP1QyTYjb6YtFs4JgRIPt9y3hnuBUEjM/4tYnmrqX+
N73AC15e3JYj/SFTQjKRW3lHNb7lS8dMIxaM/weMIZxhxL4DyoYBzOQ0pIhbFht+
Hqq72YjH3iNttPZnM00Ql08ozJapDLDgllVb/4YxClx9CFgTVHE88x/V2PrX8ki/
zzl6PqZJFmgfBWDynl8hNb8nvKIsMxPmyYriwIdw0D1MVMYxBjPduS8IgJIe2jc0
GIM3dMqA5GXkRoWo/JIUAetieMQvju+Lnvv/kdip6Fk/frqHU98xBz9shScwHArT
FGj10ugcafw03uSmC/i1gy6v1KFyne1uFr8Nqg/fnRISBeOtNoszfSxfHbdUamdo
dU4eQhVDOyBb76kGswE9Y9aBJMyIiJh0U4I2I1lA1zvI+hQSK3mieKrRg7rkvT68
F6kp7pYTJj4/+YV+tiR2nBXeWbQf0xjumfR9P4DmqyUBaAOd/Cp1d6G+MN1JuTrF
82vrjP7QTnpkyo1E4MiCYDQOE0AzZMB80lLaND8+NSPQl4ILzsAnmOV82p3k0Ril
oLXrjZjTBdUG3LeQ/OIURm2+FttCLfbBXaquvMgl84hcGHMxKrNcvkp333PYUvtg
VqGIUfu78+v/zTenhGjL+yvl4tUCDYxndPc///eLjo2BUOTz2xH4CfkudMt9KXiV
om2u6VUt9la17FxfNR0X1EF6Evh0aEZGAWtmiZf8pVimc6mdhUtCs82uEMJptJUY
V7S0rVw2HK5o5iLfMFakmyXSU+psJoSoRYv4yb51k+nzCPrqMpQ4xQnA265gyneq
nup79eU5jcDz9RbepQVtFPGpBJdlQSJTu7lr0XLf42GM6JXmJoUmo8AhldGioXJs
sYpRb40qrHGZpJFjPoad7P9KHM7IFUpCSJt/towEo/yX0ub/Q4MBIq+ftNUxrNQ7
zMZemtD6prjAO1JgYDtpYpkbtU4TBICq5pROfR8ikyZB7yZSvi88q9ypwe9WvOLV
FQJHW8gDPFyts1cOM4JCIcDbTpP8RDcpf57xhgiUn5VSO+lRDkc2s3/mdDXTWj3Q
eZZ7bd0puUETaKvlDJdIM8bpB0Z94CLqqG2cbEVKeBoCYo/oAlSHyEzu3WMEZBrW
T2C6ZqOrZzFFsG9bb7kqnhZN70sqFdjYvqsfm0H43FnLpo6CnxNGuSG+5AuHTXnj
f5H64rdQyjwG8PeqSOhLfIPUTkJtpnRuC6nemhLqPPZDRmrfp+viII/oFVF1FRmr
1cMFwCwylUD7kA8M4OWGVHaqIx/gaN7UhD4WhKdtruQdtlumGM3iNmygc5xuxMWB
5QhCMMrPEn7uBC4yhXiIs7gTnF6BhvmFPdQ7ZR4g7p6TSOosac8vnoI6D+PBsFwC
1uHEaMrl1VKHGvEgeOQvDMIp0ROJsR7ZfWEiLPlDoq8DxuvKwhK5OwLpWfoAaByh
trFbCjmbO+rCFvWVHj5V6Z4VLOwkgAvLbaCwMOjcZVqmnwqiiUF6k3j34+PkeoTH
WhuGuA0GJUaK/4wvukbtYPcrwuGLSmhK87sXWPVrHO1NXcbO9J1euQLQYZtLXVkR
Tzf2wogPRyxd/+k8xpygfShW6JsxYQe01BSmAp7re7eeyuPZ1XiEAZOUyomuKN5I
IBAYcmw8bCmtiBnazS6+K62uGgufwjlbDVRc12DoDcnLJOC42UGnq5OqYSwg3ZjN
EdMu796HTBcWQ03szZDA22aK8bTPzZtn5TGzjXvXw+Dp+IFo+mSWLjVuu50h+tdX
`pragma protect end_protected
