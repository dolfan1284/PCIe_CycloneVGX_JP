// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:33:40 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WczgUSjQTmz6+nrkMU8hqladBYv2TjO6QYKuH/83TlrDp5BZ7onQFD2ny5WdSld5
t/CDl9lduEkWE27mid1FeSZPkKKbH8vrU2YUTSANBQiMADJkI0gcynMDFl0atlL1
/cjWuq/T9EdHf3SSDZLzgEErBvVR2L8yngREEjEmjF0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
gw7rd3o7vkoe/bmRsQ4PTxfM30bd4siw60MsLVsAvFi8ev1SqIPlmjHcXZTE/FT7
oOkpnu66m6fbVI2MBHr86HKqLYLpHV8s7MaLdqW97sV+8X+/7E2vswPFEokFmSiD
jskvn53fWKmcCbJP9/KF1UuEub99paEptbh64E0EaJuK53raRsaqd12a8R0HfkWf
5ffWai4xOEA11P/+tS+Bm6p7G8b8CnMrvPOgCGHOgV12IZt0V2wyrBX6YMGVM6bG
httKr8eaKTk5x/XWN6Q6hF1+0nIq37xH3zPgf2P8efwdrhy/hSLoqL4XEC0Ij82x
xZqLtRVGOqKIRVjKQZAJQQ7ovJN8XbpKKPQ4pJ2V1+s/VRWtySVvJcTojrBjrdiv
qAI/M8J/gE9FRGDgIvRtmlYosE3yVioiHqRYph6zLQbgKfdhQFxAod+hzreWgM1E
CdYebp6oUX5mGt1KkW5D4xnEeXIKEQIDcW3H+f4FHzLriflBxmPGdDUzm+CEzWXP
fLPaYF8APRLNlkoWPU11k9UoW5NglV6wcHK/hLjcR43mY58EqYiw91q1mQT6vGEb
JYB7/Nn0cQgPdNwxkTAupU+B3kb3YRNHSooFfYqyWt9tzB5RWzJ4Z6GkHagQvc/E
SasaFS+retShR4YqFjY6zdIu5qn6l42/FddybDWjsQ6eHtHZycbaimwRdvehD6bW
8Av0xRBGvvgXKuurueGqUgLERAkR9dYcu/b64RU7IlGOsogsy1y9kLKsCm2mjFlP
U731WYwOvjEwy55H3buWwsLJXVsuJUe7YjD+njxYHDGMFMzR52bcoMHgH+cf6Ku/
KidJTWtja4gxEa1m5hYln7jmJ8MAPiaOGMqFHNx1PUIr39MrS5dEL6eM/Or4JvL5
pvE+oHlEcBnQ68U8Y0ixg6kgPaUK5fN3oDiU3cnPENV52E63yrJzae1Gr8FI2icG
g9LIyH2FxNOCckxhtz7M69QZvRoLHinKs3hwveObEil0Hpo9j7Xy01HpHDf2eM4r
W3ce2iXKGOua4yCWzjok8aGXG3CMoRckMPqPow3SaiAWk9vzr48ppEkcZpRRp12b
hbkjXqiopR4oXC5y20bTrPF4w+/LzXDUzATtZDeBVtAT7dmiVsmOxFbXuZNouZ9q
4z007PALcpJKBYad8KcS6uHOWzpKjmGplyYJCJ8D/xEKQ6vcoouOyMG2A/2ArpAh
KxOXxqxvLNK6HC9M5XPkhm2yg02gbnhQWEeExoYDzEUhxt9vINRHOqNEEGq8XdAQ
trsESbwI6qOiZZGLzRhCLYC757NfOcv+QKT/HRr3dTyX+K2VNm/agpluMCdwMIL2
YTPXqhSh39qr8uFoynEAkQTKvi68nR/nfVEZVV0nJ3nFJwmefxqu/xDXWWYmnU2S
LcmZgo+apmE2KeQXx/O4ehC84V8dj1wjI7Imxzly7fcopvo/3NmL15Gn6BUSxbXU
tlPMf7tl2+mTU+qtK0y0dyiokNpHoTkJjewhw0WrVHESBtrPC2ugE6pGhe9DZGGL
3R2FpFWCxfcoLsgU+L3EzjtVopL6V12Ixo7jJm0nm9jDChXSsNVyfiw+9ODOrPNQ
p0J9avrp0CQs9Y+tw91ANUzClvN5eHrB7v1vB6haq8BmUWjC4crrZBfaxUQNHy/Q
EUDtbAE95oHL4nvQ/C7iQIuiOxUDaBk8t3zoCgrMwuUAMfpXbYCDRdbHc9dU6jVe
5XXbGfvW1pP4MZ0ZIIwvIz865FQKoe2nm6qF1aG1bWaZUitP2z/49b7Ruc7icagg
nPh1jYhU3CHiCj7yzMv5VtTYNv5MsUGk+0rRGRnTKQCXpQXskn2NEzWqiBoR2447
MYX4goXPv0943XVEA359c2bwM/d9w0o5D/70rHSlWsc9U1Al4jj/GWDFBp/oz/U8
2MaVjMRCmx7DW9dBiBWsrE2SqlXeN/hs0vUrJ2zq2CkRO9VdbSlFXpJ3KQnHLtSC
IuQTLDPQplLtAnX+hvG0Pl/m4DBLnKTr2yPIzoaTYiHifcg1CgZs0Y+OBCwJyxVQ
86zVfCqF5NuklfqAGF42qR00QFcr08rYd09UTrQ0koPBw5I0Wod2cDGfl6lwz56C
PsrfqzwBWwgGKJMndnXqkjiHzKIDkJYzv4pTq0aECiX56OGHqnhLSclUqxGvRMsH
wOtmQHz0V7Mj7Ck8lwNsoC6b1CWKr2mKh2TuznvEzv4/ArzrBEWMpz5u6LztAeek
wjuK77cqwYSLFEPi82mvhmM8OiF0GtTxBJg/zct1jKH8MXXi+giDXNCz84wHu9PR
tVYjR29zbBH1X/8xVCf1zQtYTN+tXMqJKTUQ6XsxrGpUA20/yPOucgmvUW9LGEWx
2TUpHiS0Xangdua9Us1xdMfKTCdxcc5lgq+iC6u6W+K+/cf1IF2VmMvXTal+mzhJ
/8Zdz0yNUyX+jsv0dot1dOb6qRw5bAjArXTQxsaOohezRRBxGnuLdOLPE3SoIccp
k6P/ntTdGPDJcdlnUrL4XmcgQNjkhOtBzvAgS4ua/NkAj2lNV+wZUG+/xdpDDDJW
ugmS8YuyI2BZbwlEOW+81Gw5eU4lZNJokEuoKnC9bt4GWoq2PudjUkTKJieiaTFu
3bavltyKtafqdVScYqdrxvHbuUY0HfqlvG8KDx9zcsqdG6AADQ7p+uSwq6o6alSj
Fs/vQScwAlgTJqjtmq6wPc0gCP3rMw/LLNFWzHX+lG3NvUMzosQ/kCELMm/VlnNx
BO/ZBXEwWg+VtB2zFaZLKKAq99cjQ/Hlep075b2Ut4uhyrqjQZ6XWVBgYSogr2t6
AS+ctZfNVnm7nlu5BSoXcbNZbMgwJNdzgTkh8VTZiSHf17jqvZhxrL8FBObkHjX1
P4tZn7tJ4Z1HEb8cBXnTgrkAHN/Kjl5vd0mJyC8dzKRoG1k5xo4rQHZ45twH3wiY
ZK/7XW0RDoMl6nZRVEq80/s9PgHh/ngDa4RXzsNE2InLlaEH5xMWtaQOMu/Gm0aG
zitrp0/yF59MqczcJpjlPyKaLPeqQ+OpYIPDuWNU5NOlaTV2Vo2gyGmthb0pyR6X
KvevmEf6ZQYlU4vAgf3xhvohnHrlvhh3neQpQtPzRM1cBbXo9GeAcGWzdtXKg+gE
2GGuOZ4ezvLDJlgxmtLTYkluS7edZTx69nhtdR5Zf79FipTLDGGavgwYIJMJd6/F
aIJKFpWl8TLgGFClRPJABS9bbR5KvhbfPwHWjzu0QDpXtazIMbnM0ZqHurgYGDgb
nimpz5+zxEE3H/e1j9sQim5pN3B+/dO0g0H7EvdPsSEt96nNPwZ1ueNTIAOXpma1
ezvNZtD2FK8QnFrrPeiaLlMK2CZnWpnOoAMfpQ6VvaDWEnhMcKrIqycX/ZGEl1Ta
KRCBFBtmis3UP41vaTeb+W7vyIbRXvv6i9uxxgu92bl1ATFDyn/ytXhjYNDBHShL
eSuUdGyK3UgeoQpwy5P/32MfKXjVi9z8bx+j+3pQtARKYDwESpKMr4UXM/PVimxI
/EZ4w2IpQV3GD/GInAiv41LtFrKCbgSpdHqs7A4dQLrmgfXXcb4w4z0PZzQs6Mkb
sLepqZm5K8DVS4OkLWL4tMcps1hYcsddAAjmBvWV2vqxjAAMzos4+SakVuKgJ7m5
kTI5DUw1kOBk5ytmB6rdcwznxg9atonBxNN+gz3CZU8rFC3Qg9lGabZ58wMmnVdn
8D5zh1CqPv01upPjSR39zYInRl4GDMO0EoiylJf2VlQp5q7AMjDPtjvbjS5U9XLW
5LYIXPeO+YtuDwD3onoCKTyqLnwEFnaRObEwwpNEbjZJQk4IulDZAkiWAb+gFsqJ
lTPNur9Z3j9FgEp1hohwFqnjqI1ywNhg2h841zwCuZOxNAt+WXOKQdwCzSr90jBw
/u53KFhna9yQXLmGNWLDfMOUUDFpVEvfLrSIeJv7/XZtlLV4dlTjwpCefmW22AkU
FH01nuCMCM9L2CV6RmHDNL5m3yXQpr2WV/AVSh2oUMwr/NKHdali7BOvUgn69+fC
cRFdp29VPrVJypre7zq+lw==
`pragma protect end_protected
