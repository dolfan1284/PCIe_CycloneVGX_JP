// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:57 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GPn7fJtoRkSgyRLSgHtVrlu0GOwK+3JUWV4pHfZm8YYk0mKRcJbePLR4ThpRXglD
S+VOPRNpoGRpEIJD57Y7BJz0DzTYUgNzAWt4RKIvwf/K7PdALbPEgTpasmzesrUT
VrmnP9e+Ox2OCtGcLKwxjdd07TB1Y3gwqLkAt3FziaI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
9IDejINyMNlnBaPNezgYTM9nufVaC1WEP6uA7XA/UWgquxTOqIiy1EGriiBz5QT6
6l0696DLuEHRttzRMEOYy6m8Yxj8yDzWKIQXBlJi8pR6w3lcqzZ/LcZ6U0FH6QNN
nlEotmMviANRaS0ZTjYpc5O7Ej7e7znmQ1XvfqIguNWj4EXesMIGOexHSiIkgrKA
TiHEUwhdrtn1E37hwzVDVfBOx7SWzKXwl7vm/pennloe997Qhqpxr4WPR/rW3MI5
qu5G2UYN2oWGlU7TcGnMfZueTeGkB2QF8JzLGzLEzly9LexEkkmGNR1ptjuPF97i
HQWjIblWhMts1VRzouQbDS+CMuId66Rx+r5jIGJMRhWK2Q9teNTDh9/xmRCpXJmz
rzNJ4cdb+nB5cmm2i5RaB+6urd3pisFOHcyIGHOAN097RJ3RS+4H8cQkrL7DjkNa
eBfjXL3+5WYCbkjjxEoMWSyjvToPPDPPWmcn529Cko8PD5RGeYyNuz7O1vHQ9gQc
ZpBQ4JVsFmwQEnQG7A5FfcXd1xP3X9tNNsWdRd5JDcg/qPvVe7IQHLS9ySdbIcaR
HY5aB6L9Y8QS/B1VkAn1pbIYJYrBQl3E0A0vQVP5nqmyHOtySVi4H2Zdo5TDrZSR
HEH77/9Yz9vNzSf9qLBOh0MiYjjPROVnLMGnNmEQyqJSFHbnX930sb36lY8rC49U
yKNovT2ilYUn0Rpvd6J29ZUOFNBGcaZiit/gBq7AZom4kQT9r3V/CEdHs3lzW+0h
IFnyj8A9wBIvzPxV0TpYSenlQUOeeNiIBW5nmLholptqnAhHOlzo65yhFsFktq04
Fe2wyMpEj/iJh5gLbr39bURDM9QMF9NfCwwSZJe4yTVTvLKEz5O+TfnWoKZ+I+CQ
WAihij2KipCNP0s3dSwVUSs4Az87rat63J/YEgMjBl0SOKsPj73bW6lWoI35fUY8
rQ9cCDVs+bd+OkGaWFC8tZoXEQoweUvQwt/b+4BOyZTCvFf2YND6UrRb0m4GKN35
JQvnfwJunIEC6bO6GMMY87bixNRQzOYIgXMEDqlOkhx1/CRZIuK0umqWTz/M89xd
yOQd0xA76RdJIHg8yZ6DfigOYJV8lGdTSqEM0PyJ2JmIvO/y1zG6iNo7C0hm+6W2
JX5uEwmDhFATm9Oo26E1LB7GR2qHiObk62r6vYfMM2kcEEh5CqAc2G1mO0bfMWSN
67uawDfzapiYHwyfGljQZ/D2JUDb7T2jr+ovhBd4vaQuOYLreL2zcqQ4JxHmtq3K
WI4BcGgRfuk9XBpgx7ICQPzBNmYZoWnzaaI8iODxNteuiZrbDmi9fP3ECsO4X3iQ
iDZu+iVbMNzuPbjEMmhAN8vDyBvNKHaoK0jpP+yFIUsUVuvaeqX37ok+hfoQDqDv
6CQ5wx/sYAbet4InUpHCRy749OX6Nugw/183V0UtfhKcHEEjRkK51Ty8WuaOvDFG
VfwWBwn1kl9k9Oi3f2t2Z0XmB1KJl/Os9DAKcVdPx6vmw2rgXghmhx3eRRlA2oDo
yK5zRDn32HdfXFwBoy69/QI9WpYOpZnlz7tgYIioB9vHMxojnlNZ2JVhmrxxfJYq
Ga4oPFyaFpflFr+CnjtB7NAzcBslXha+BwLcsxfkh+kgEU5l5eITliIet+TlX5Dq
Nnq+J9I0z/xssHf/y9rH1fXWF+2ucv393gse6RpL04EbYOS4dgXNEsuldNgSjPyy
VSAGK8dofobXlpumUBjjCxwqVV5GsSzh7BKYCi5G8KsVw+T1VzsjWQxqsPI6yexM
RdVi1N0FKLJZPzOSF1+XIkJomFnZa6b8jFELxy3MLP7Md7snSYtCezha8ap7h4UK
G/MuxWjVipyYdPNZ82r2pkS3tSg4FhL0/5akU4WEJSR98g1E8JJJ5eqIJ47rMJgp
mTSh+XLmgQNm21pjIu11A9GA/M3RHKXCNOtF2nYkR1HHKrvy/0GlJSOHQz5oR40k
qviz6UrCf1OMrxQMbsZYJZ4ISRyY1zVW81Ac1MaLxBqTHQU1DzzaqVzjLNscAURt
NkmuNamw6S5mGXJt0wyDOyQS/O6MEZuT9lnwQm1rCzBjs5exR5xOuNUFeZm+6hnI
iRkFf88RajMS68FPxhKtoaXQKAzALSPeimvwRrVc1HCZ5CrAxZKSmgV/0tvFy0+X
+WZa1L46EXWrg7Du/eE0FL66qg15TMrA/K4nteKD/VZZIYO+qkiBm7psVHv7oKpT
FOFLIt4Z8x0eiRWLs9MRrT+PI1kPqi+WZO+KizJV58xOB24qZJwaJuo+Tm0PWMaF
HA1pTpT5NK/P+fv9c65D2PdgpRrX1PcSsp4aPjesNeQQGMiLJZLAyQpzHQuPfzDj
HxDd0Wn5zSm1mx1CO5+AZmxGbskI5rbhPwfTqFlFYPTHmjoclN2lkZPJgjrx2izy
AxZZkbW/dF3i+DCQBfNg6SzPoHkvBucv+YOA2Suu52D8p6I+00eOLcG01yPG4lPV
ufLhvEc31Zj/kxm2UpPuuliZ9PHZv0ZOiWdaEZtBw7vj+O+4nIDuImYpDsBOHid6
DmIOIZjHIVuyvcRCtaQSRGoWKPHdyf8YW3sFUZTjQcZkFe2CDjvdXVGzPLsjAd5p
foUSJggtjfTMzVTNkVq3dQdhV1nsgHTxxRshaphFSfuxoAs2jSO1edvEblKqgUVR
7gJrdE0hlJALvYk0EEpxLruK+O+TjDkzf07qZ2eLqn0aYp+tsO2rWyHY0M0LpdwE
eYQLkCyfg0Sl6zWHNcHRTZsTFNgFSvHC/6IwmWylrqrly8rHiPCN9wv591El6ToG
T1rpdwGEQHW/gfAYXH98pmqwnM5nYOnjYk50q6b4YAo80OO0lZTEg5jGA42FE+kt
XFlduCvhw9tyJF/5wWw9/0PPkHS4Gb0erH+4AMLGHwykVYT/QUUQX4Nap62YsSbJ
pzo+ElKdANQVRlUNiSNxz2H+YFO+CfHq6ZFZPEs6MjevWls27eKxRYjhWnnTWqY8
A0qMpwxOOFN1/n/KMu2oktvLnSJa2cf6FfAFyH1R6XKLycYGu1sEMAc6492eACYn
oBiir7ZBzhlGbPeInKHQAwQAyr4lF7Fzs6FhuqMlsMrG+B9PNafYXQYwN5v8LRHE
xfj6DLj+jeOc5RzkSpr4fCKMDaPUsr2C7RX5xg+LQ2lIj5TBPjvst3eVhvCnMvTy
cgw8qgu86bjWxXArNjx5+2mXwUJ4Di6Se/D+eVefYRrDy/lNqpljJd43BerG+0pR
XrIiMZWRujYWHACjJhJcm3yWu10Bjdm8nq+SQjNXnS14enJb8XVOEGeCWMaovfMh
PK///8dLZK1KLIbg22ZEY2apUzTzMtzSuN9CbYHp+iP4b2m1I5gI42xz8ykcHRls
P69sVl2su2/ymxT1ffaDdtxFsNU+HwB5gfuc1M6iyO4kWKDgdmrffpbpq+BtpJla
WpOeTkuN+hBB+MxJOf9qd4hhR+0ELfrcMVJCiRychlWwJD4ziBWRi3Ws18Cgjyp0
k7/qBcaOXo/oA87AQfTOxqy72L/nLwzzQztJ9lNc3FdKFqaSeIdf6gZo8vjS6REC
k4q7zNdAud95l9Gykb6w+HAjoGvPcKsh83i4EiKO1SPIy6N7drwEP1nI/nEEiosG
IfCXs+sJHXJs93dXCvZVMmnrnwVbeEin2pnA96wvN7IAQXENieZHIVpd2ZwB2JD9
bJfFEbuU59jl1Ky+k0usaKP6Z258uE559RqWvbPhBzzzVNdcK9ovYW0WJgmCkO+Z
UzZDAIlF/2FzDgnMnGQYwqQRhBqVs8NxKvxwto4GHVMRzaBYHO+U5u+QBHnHbu6I
1jQS9n6pT0di7NOae1y2nQncKy4q+RLTs/Qx8yhKNJQIsJLbLB69nAAlIuMhi/cT
nG6vfE5lIgFi8D3/hus+WvkgKwuYv2O+B5gZc2dFbV0id4vSRQhKP+si7cPKnXTR
vWZ3bZ1iOPDG3vg0tehhwIJPSyZtAwPMZobQUfTVRJFZ0etBS3JkcCqNEIPhDAhl
Xdn0g43yJHM9zTKXyXtHYA9DfHjui03yF9m7LfGLzkrp5RDUfTyezJpn7jtu0Mtf
rZX3j2GffwH4PwQ0mv0J3/mzxhPoUIegznGHQd2nwmevC4Ee77Dt/13IA7YoRGzY
tDkUx4PCHerOYeFj3c9zNnc/iOCvgNuVxG1M+9zNy+R+z2TpBo70HT09D7kZC/CY
Ays9tXAkm3+esapP0KmuNvAR5L6VxZYJ6SWhN0iLeMe7E1/WCJLun1NfIc4J5Ujy
Q85b9HNtEQUt25ne6VCQPhrMSsKnCC7ppvi5mcOITiAaIdrK0IcPTDeU5O6YYhe1
yusvQZTmrDyWTxLKMNJYNwoHtfGcYz+CJvD6QHsQbq0YfHrm9IhkRHgIwIpCQJ7u
hh8owucciO8EOiq9r1tDgkbKTBk88Z3omJPNA8x7aSBCOay97LtxyPLEjDcHK8mr
DqBK/7uDWnQXfPvFRVsRYyI9kToCYc5BlLulGuubZ/RRmmpPVAQedwsBLD/VLz4P
pDQF4/rs37Av59YNcc+wqNxBFIQ0AcwLfyursMubtUlCYTGBAnoFWrXW1kGsjAS2
6tfw75VDdXloQDBOgpvpICMQbYgXjrBoRLO6G569L4jhehWKNR8hcVSF6jlbQmaY
rU9Gz+kautvAz6Wp9+AnB+7mPq8SGqAcSZZQSnc/qg9pGgEZ8+9uFhtACvUTm4N6
VTEoUNR8yukamagNLLdS+64WLxaOWJN9vB37Or8TuTbN/wkvp5NVrzahYYdyQBYn
6T5dqOkOqu39wvq1SnAHMbPprgkqP7rVmnjajWTdcZZ7h5kQgW8Hgbr9sG16CwXI
tAPfkweH6r9zNd13tB7Ja8sjxOFzFjrETltX7Jx0igv8XrXmHKKZ0VxcUahTr58Y
DVSisumOqsoTnafYgTPpicxMvNBDRGyKV+782m6s4PPBOZTvaAqxq11KAaegBQQI
0uEb4Kvm0DIiWlu2oP5532b+Wn+r1FCKBBtUN1mWmkmufo8etjv5Givoh/YMJZhj
UEzFFAg7wZIZmYi55DR45NIR+OuQ98qrkhDGN2Uo3oNxAuPgS+4R5VrOMB3MFAfg
qnw61Yn9Ngs211hsJEo9AhY8BqsdzsBEc0QyO+gNvWWbTumObbVzcv0RmiYMZ5DK
jgVOplvLjT/ljQZpGBM2x+wMeW5EZFcTCIoi6E+6xRDjvWhovyquKkm7ocgJgqPH
c3eYxnhuBsMH5MWzpH9RZ8KBT9gp3I5goOoVE4sRRIcgvV19hsD1g7INn1MgV6df
TW5eKiw1ge8zjIRUGSFqog9OmSjhmZpmN6rTFG91HWBWUectccecAhnG8L+MeI6b
zz6QcP26Y5hwNwrWBgoXKb/qWYrbY+Ll7nKXlQ9zkt/GQ+nNwfi0cHR1PSmNMzMr
mEDfgSsuPk2XaVNN8oh8hoK6xHKHDVrXPrZ6UXN63R3qLD6fZhFWdqC1N8FgTEAz
Acr1Eq0TUQMwCXEDcggTD/fCMeWbc09KXOhiXhkYTQdDLy+RkACNCDhC8LCORVW6
NsU9pHiNDRe2FnI3w45ZhXSentepeUGC7D6pINDL0pI3vWKLj5j0vAfRThHvDjT+
jta1jS7eoBwHRmMmiOqKCQj3MOSOv2X9mZLMl8adki0Xf2WXfmCPv6wzp4SV4LEA
CacMXzFnsw5fXMhPGrS3aQRN6Y989BthIQV7k9hgbxSal9IpL+JdIWvffm9ZqFal
jVTmi/aQMz5mClqVwRibgnNX8+/DRFTOO5V2mLdF7FNNCzOKioQ8Uw+8SQDdxOlF
18vLJXK9qJrlpLcpnsgOBYGKfY9XXzhW1dK1wCxYHHmuwFK3hyHx7n5hbKqDhl3Y
04dA+pxoLgIaumdwQ+frGs1tO7oEYMCcQzYGFqnVEl082321X0y5xMItIVOHWjWR
POoHd8ysJeVV9lCC5YwVxEWqPTPd8Za5hDcdtCAtDKMVXK66t9EyKChP3XJnhXEj
NWtrvpZoAVvL2EhvmOdi1i0Ry0qIMdo3pwsSH3xVA/pQ36WX/MJqFuRhgGrnb0Zt
DF3KHeV2pToe54c59EPSyr8Dw9xkYOCGZomdWFQObQOtLlqpKDwT2o1Gw/QenbyJ
iX5R8sDJI6vNh5bTlmw6S59RtuQpBlzri4JN0zdurK/tc0EdzA7s1cgn3w02MHQJ
zfmTECyHMQPaZ4vvt8yVTydphTlF4BXRayppntnPJA7oNLco4BCBOI/evQc2gEYG
Qow4Azo1TgAx3Nwu0um+T1+Wwnw29f14DGaEl2XfYYldlyYJRbU/xwRoJ0NBjfFE
/VrJXn9qYdVJ8U/JsuFHgycAbDoWnpEpBbNz3aj4CDfSmC9MmFXCdEAbtgmANWLO
l5oPtLDUNWUcbF7Xf+Y8FxeDQEKpGP4L7IKYTHy0bZZAD/7OuzldnbV05xZhguEv
ZQLzUXPKScEQ7UlfuLQg99ihYH6F46PwGbGBpQZhrYulHDWhhqBQSIcDXGUgBLoS
i+kdEwItUlcAvCfLh8enP6luGAambEktN0aY3+Gtnkv/Itbg2ZsxZt54SDpXONh0
/4Dy59J/BO9cJNy0IK+6aHWAkfii0LC7+7Om6wncJ1hJ3O8zFlEEZddwQXCyfczA
9lmuX/rAmphbQPEvG/qbX2MUiHXEqBhdbfYbMTwFGWj1KCGPwMYqF3RUVh6QvoG0
bOSmRSEGMQ10+emX+Ds4uoEVJuohDhhq53ZNagundqtp60XXo9dTn5YqXANxIdw7
KB9u+sBNhnkdfEbEX/GiCXRolW8vJV6rnPYAVxkx0YYLk4ZguPCjVmNjNuE2kGcQ
jk0WyONcdRvHw7MybTiOqiYVdTHc5VyHE+HCHCX+yNc5lVgl88IeVnuXXZBPOoNu
cVlh9kK0HwIOc89vnutZ68d+qvqF7ory/1uHgoDqHIBEtvYvu5JxmAMwNtlAODuR
2VDNeYU4+27QEVZyc2fR85Mtys2U14FKGTJuHcxpSmaRvBGuTWpARmcK6pFvZHjh
CwedK04mUNvBUhK0XMWBcaYnvHYQR9p9/St9rFzlKTnNCmjIS76eEp45RvwGRUsP
C6mtOt1a7PoWf4167yc2vEinpAp2hrvtQ/iQlDR5AkXI07kZx2BfAjDyHPSKtBY1
OwUoQHmpMGoKA09+vLgg6RMkO1I/pZ+GsRvEve2Xv0csinWa2vV5yLWRK/PHOYsK
p7kEC7Rk7IFjUFLQsj6XHBFyVJPmtxQGsz6kdIl4R00u2avbH8MamLfnIIYc1r4K
wGT1mZtgwvMAfqfR0TtyD7FwJLAv/lMWkIg7lfU/ZfA/bnDv4n1V7HdIg32Zh4zH
YN0en80W9Zsa0JWhP3F5KHu8xAM/USJMfo5l5jpFtJU=
`pragma protect end_protected
