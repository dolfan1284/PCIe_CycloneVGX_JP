// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:01 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BPXBtOmyDjeiU2yiI1ihKk0wSIPKn0TbfWu5QOEhcvUj4tpFPmNSjcb9fCgAX6yf
g3XWvjTHORHdSclWNNqPRozxuEyLbzsfO7MeoEFCtMyLmLdlfSim4kK7bjqeI4z2
1y1f2VVXWuM4cVMfl0dy8r/mm/kWvNaY6tXbx42vCrE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
c4tUDJYjAn2PPiypTctKpgedN+0n9/xJBdxYTTznbTC7rNdhiPYpgNmgNEHFQ6LX
LkaIYOpiVl4VKPXTz4K2ILDRi2pfvuk8UgO2Iqv79xGMr0lWNefa8Sofog4inRmo
L/Zg3W9bdQeiLdtKQG381d10oVTIGdKzDXwE7FdsLCGNNzNq0lV7C9H3PwrU1Cz1
jQvmtlbHpbMmiYfSISZCX1gaQAGDfmkX0wcCh8zL081dGGMJcYUjy1ZDLbvnFcG9
lNrSaWvGGmhMnveXDUuwe1P72hnfMgTAuU4fhCaRJGJgqcOWbN84KGf5VA41L8kp
TcApRbJp+nLH1MVdOa4mURZqy4bytffydk+5D46i/POG2V2CwzVPcHsd+mjpjiL3
CREhxyCFCjVvqftCKntFndoHOHWNF9IYOpL+ADAA4EtKKVCrBUogamP+tKdx+IdC
VjKmmCt5nPdjheydTu8bUyTBvjQNpegz7ztG2+odsmr0eS9pepvry+KhYM3anqBL
sDuuktty1ozmUT+cQYvFCuuifMvLgLjsJJw/bl9OhE8ElHCaZWer0RHZbSNw2N/y
/AjDvAgCEM1MmucS+JF+zEpWlDV58ZDE/aKvZu56ueFA4iQiBuVKryz8kNHpuMOB
1p542gtjQzkQB/2yVvfOuojHGAlKod+GmO3wpgMxhagI9ug85nfvpSulgWlesk4e
KdDn60Hy8qUA3S0vHADj8aeH5YaBlFyOWASY6ABQKEmCmXrT/hxpLKGUHCpWiKu1
l9zAYJn4BpLP6+dNpXbidPOnq41CRpCcNV8UaeDp8qgxitImmfcAKVfPiWKS+CGn
b+B+TB2cfvJjGmDnZNScNLuhSdpjoVa06SXQplImpzAWplsfYskQVeGnSZAZECx6
AwJ9KooeK4RweX29dsU1UmdOyaHKsITEtRFmFpi/ZHvjTqSyK06px2DyvmRqezJQ
CaoJ+olPBTDu9R+h0QhdXdwajCKfBkZJE/xdG2MUFrhwQLWPBBqKr0aq5NYtcwUn
Zh5jpVmw8WjeK6puDSe7TsWOCtX2G0FGk1wNMd3Wvd6ZFcmctXdGM3lhyVezv+na
ehdLuoRzSva9WXhjWtRjSeHuUwa/8XxPuxR6fs8YB61KA67RX2fqtU6mkbQK1kxV
RZeq+XNriFUX9GPOMguAimFe1rCQQpXWKAq0TnjpH6UhyZiSJnvfzlQiTavS5zzV
3+X8P3Hy1h1At88N5axGVWE/HeGE/X4iKYtAn45JgSd4O00XhDrQdDipKb7hUN06
Kb4MvNVlCWJh/EmcHIgXyPwBFQkOtU3u3KSYwJzIzJXPTFIPcDbVfaGAanOPP8Y7
9i6VfR59K8XIWrgunT0y+C6uw7xCGb8xmjj4RsyI7AFaeleka7kLR19kM9iAf3N4
otW7SF26M5+98/Dc09Ja1a8EfNo+p//58v/jJNQ5Be56PZaDwrnXq5xICWOMgv7g
xVx5Jq0GUahu2sr+fDXcrxoem5ZdrecwFZbpmCyQ9jZhzmZBcLdRYg3iPVLdI75f
nZfne3LqpDPlnVZyB+PYAlgjCCcctdFbOwWi1fWWqmLDvUMEGmWmcVhFBz++QGXJ
ULG/uP2tgUohYkAJdqGzcRuCQUU6mjvhbL1b03mlXVgSRUFU3Qzlb1SDTS2tAAgO
MJRTNftDTF+d9CYclfLl0DXLwKcKyd0tBIBzv5KseRbat0/M1VCTEGWxHCFqwrfd
m6H2RzApCdAK8sa1I1wzIOtPjxqmoqAfO0LmmkKlDEVrOa2X+I3y3kkbex3G6N9F
o9vCKcDK+yUdop1/gOnvL7U3BR3UpfwltftCGWiSeyI4SF6SjVi/VTQE6qqLxGZG
IpEt5zwi3eyu8ki6azU+Q0ycmAEqLA+LeUcR9lvEqG5KdNY3GXEwx6Nns3oommpl
EsrtefblzhSK73USbVq7GtDa5I2z48ZGhRSayz83mZUFB4cllBEjjy6M2bjfPNVW
+nXvfLUB1GTLD/lQNvVtM2IHUi1jRxZeR4e6Skvbg/eVsZDNAhKgzj+m+UKYMpFP
WuJNYuBeQfikJBAIkIsEAxTSoUQUcZFlDHFDpKdcVHEm70U+NyopC8aRsPyeqTsE
Alm2fG8UwgakwDXoXM1Bcr9G5kjBA90b43AfBcTH9S8q8r0jPTi8iMTDidDSYbb0
PTEMOARZq+X5Z3e2jD01OTBkjzrtJ4YMv8eSBLeIyZ/RgMfAzFA6ASCqI2hu+Hy/
5wtGTgTFe87M/m2aAJpxpxF5QxiNKszebJSCXmp+0YHH+ztrBBn/VEZmpZu/OXH+
uTLaE72Dp+5SmjO06XT71AQxN0wPiihdhWIjsZfyfct8HvQu7oi2tjXDErFQduJO
XBo+lS8xZzJ63J0wHNC7PFGyuy26glvJFQAWkHa0cKhCG4sy1pcrkJxtFnq9tM5i
aOzSpalhQhunZ9tqgYfGeNKrGyxWNa6qKFdjMh+UYsUYnPYVAo031cJBi/0xvBhT
7g8fGQ4Ur8x+bQBq7uCCK8U46ET62zD7mf3YB2zCjPJqc5v5S0D5Q/gml9PEYzQL
YWXvSlEr3WJxgbxOG2YDmYlH4dvCgKEMnqQQjLQ1rqm2Ayk9oQJAY46Om8o6mQgv
/zUZapCOvc9/V8cQTemKCDea7V40tLr/1ritn6hvIbg23ACQL8ESZG3h0PSiTIMS
m5/YwrdCMrKT/ugY1b3OyYQK5WI6FnVvNtSFihH3EHkahzFBpxUcolmJGre1reaG
M8Yr+DDBL3fcMW6a+Ctx2uKKZfbCLlnbS+AXL1s26UtBhnP5Njq9vhIsEgJmFN3+
FhVWwGeO1Dp3iKXFwNPhC/n2cCE+rNmyuwzMf9nk11irVivS0i9pGGupjj8l5Y4f
rHS6/SQAA61mv2qJEfswKovQsEuQ4e/h0AJy8j57hCkMrFQnrZjM0nF131B9JHxD
32ZSUbfXOPTkVMapWzcl2adoC8zUvtB0WEtEhwHFBn4Z/SK3sVtnWZxI9NuwllqY
5+SqeoMJnbbS3GQKxh/1TCrJQ6l32nGHXzq+i257sImdF0T2jXO0QegRoNw9BJxU
fPfmRiWD7n/d4eMKmn3JstMIuiggQMs5NMdimTNHViD0BeZzs4sH2C5gJF2YrK30
rXcJDGjiLNfSKgnwjmtB685eUQTuDWnpYWiCqiYsdEKrWUh2zVE55eGu3QbWr4Q3
s+wzOSzoZMzI53n+3QWwzFpgehxthmx/t/2RPGxmD5ROfjjCZWklIaCQ5khwlQUL
jKVdVjcGrUIhIoe2FBYorj7WFL4egnT6NDtpVvew3fyofMQbhZAhc4iJYUb5Js/5
QYw0lzkFA1r7LZRl9hBk4CHmInNJ8zCSZ64I0Np3p1KU0dPHUUikA79DjDcKi3ga
V1pHrD0wdZArWeOO/pOasrZ2FRmKUxjgeQLstSGuZUCb/AlRc0uJGaEYiM3k8qzb
b8NS11bFIKQ0AganZAENrnzAxROuUUqSbzbUvhIRvWV5Q15MYkWvGl+f8RPFsuX+
+U0ACWpBgrie2oPFz5nojcvN/PGs9tQ7jyr0kTgQp0VIHsBT35jqI30418ripwA6
sJSg9D/cKZhWcrmSwrh2mSyG2ZRwIF9ccb+v+1MnR+JZdlpaKWzyRIg6n3e+eh1H
uyAheHMnRioarybFiag3zDTaO8O0yD4Papt5y6phYhqylDtdtVAHpOFEFAT9gBzJ
g0g5jZGWBUAudUuA5N7ScJZynvN9556C2d1yXHDNeLDtpfQIvCZk2Ijzfrx7rULv
+gXz41z0ZPM3LhgCEO8su7PeIS4lF02HCK39EKH8+o8TIv5o2f4n+j44APlePugs
WMQIdOnXNdyN9af9e8zAjDU6Gzj8+iPrX4t1sGiDZVudqQzmh6w1ib+f9q1JPCjM
ySpKY9iIxsj7pD51xjHOOKMEtq9KIMY12ckyTuwQl6gfPsCnv/kJRIyPKyxLA8CW
AWXYyuzm1X29kgvmhdJOF2D4TJ6JVnCjjAJkvWIuqTh980ElXeexi5hTNs2zBdDW
agCRSGtyRB0VCi03+X3E+2pIUK4yev8R2dIGY94KaSYLHDSMSHRhuF6VXBNqB7Vc
tRD7C1RRr8TU0Ikbu7ddlRk6q6Eby8KEPgrIiO2qjSNt4Xkm+mZIzXlNrNROSpke
ZeGplRt1z+TC6PFiDx9UbwbiG1XXMl64tFtz0dyGRWjZaN4i8ADERqZGRiJimQA/
87EVUS6sIkh+Fco7iTEYz6j4AcwF1foBghZQOGJU2dcTANDK85Phc28W2ilY7tqw
ZfSwRV+mWQldkgrDy8NnlEnXjcgkDjJAV4CKoAsB4a0GnynJY/QbsFnZHa33hlI8
/D9QqTZtxbynNVivrjXHFSiMEcF/zpBYZp1R7iSJEdbgH9Yi8Ljyt7IDPSNbDzLk
3dbnl+l91TcPn9FOp3+fsH5YAUmON7VjQY0Ss0zjxaEt0rvhFazzcfiB8X1CkMXU
jdK2lccWwjL0vcyzpgEPrpJrv0Nw1PahwJ6MNkZ8X4OrblqFBo4jzLnsbrHfjg5I
/OXYwZ3GODDa/+hMo+YFdiUbGC69c5bsS2NcA7Qj5CMUhTacIhqZ2oBJXGZ+7psX
1l5ZKUpOx4NAUzYxb8bxHxRzi7vcvxN52m0eh3iy5mBviUFb5ZbACcaUaSWgZpEr
Ks2fdAx9TZ9KhxeD3PdsbWDruCbdr3fYKeGK7zCO36py/xqlbx2P1Cjfoap10sUy
weMalBp3AZmZbJe1Wre3Qs0diroMVzy5xTzGPuyCb7MahLocPNm9UodsAchNf4Kd
RmpYKDitVcM5R0OgwrlKgpkLBW1izPasMxNoMjl7HS/xhsDofSTyEXsHo55XdRq0
9nO2ZcI6pzkeLcGUJWwDSlPvQLwf3bcZ/A57XD0PdG2l5QsnwDF9EVlNayU5d9R3
ejqFgFrp/KwHSbBEgsvqTqTliCv1xXqyxXdeBEPwa31OFHraoio/I1UfL+IXJYBR
YOk4Yu2l2xYomZ5Fec1ogjzoML/mbo7UwM25jSivZ9QWu/YxgzwnXXRu3KVR9VKC
NF5OEa58t/dDTNbL3svuifpB6YW8rjTCaI4PNE2kqJ2ENQADPlbM6KrngYOg87mV
n9Mm+gZCQyTgWwpxY+HOvQ75T/ny6LAXtmxSkLceyFVnqVzNpGzyh2JmrOiQzJgM
ELOf/ayUe61l0gBbAJfgjDDXPoLgr5NnmrL7wsX4pMXJOprW42MqhEJ6Qrv93AEY
a3z9XuA+8KOLlL0YZNS1xQ2YFjdNgr/2mMAQ22K5Dflwq59Ur8aJ+mgBfbx9w5KP
oV9WIvmJvicmcm5+JeEcVZNc84tBWEnZULaiu2WqnSMaSBXpG1zGUvVX+0fvfEmj
S58vQMOS3+zbwG7VXs00FhcVJ7ClID32nzS9DSuACfano1Xm6L02QMeVGHPqRYuC
SLit3a1tYkkQzEfLrZ1x4eMp2PtD5YEGXZGoTHSAfU1sI324/frGDECXMgREX4+x
LF44uX0ORi2PPJAjOiv/It2nm2Bj9VZXZd3HN1h4awmbz6XiEZZz1wCxPEJtsHGK
FMiLEhkOyTr7mmdwxfkHZ52iEHxA+bCtDoejle5OMdht3wcUaChV4txGJ3DWZlOz
HwNKsCQLNS4TcFuGlD82+KdRTW/tJix2tyj4O/+xoVnHpe6QwX1iFJKCl40ku5G2
7Ly9ekMI+rZS4A0T2XohjTSqEoYsfw3ShVWsKFZpGXEmlhseXJlzI25qL2HmTt/s
Qsjd4X6enjIqFoyzF9ip4vcB6EcaoWcIGdjoCUvGscMMbRMSAetksT72cxjJncKg
M2y0l74nfYuFKp8asZvNTayN5bdkvMyHMdIQDNk+H4RtovEKVHMLpUYIg38GHu5A
XOarxdJk4U06/OMOxrp04R4uVqsz4Ps4guiEQIkPrTeKgCqKcLYCNPJNOA/hQg0w
prbQIe5mTqJgXqeoMDitPAGThBp8K/7Uhl/Q7KGigcUY4fdphsVANHtIvhf0w54a
y9u0zXe3zpQ3nVt7tDCwcudP8yMRs6HrD5JV/5etAbMb5DMgUY/lGMF/8KySlKSl
XlLHd1uA5AiAojiIXSuJTaBGO2WNpwQ9G6SC9xVgLhLaEQsIIrc8Rnrb1bm14uxp
K51RgeOVucFhrHOcAeo5CbgJeJp+qv8TzDCFnnYu+VB3owdCHdNrl1KRVh2Em6sc
oAW+ii3MOp5K/i1RSEqf++RtwaHticAsaJ9zaxWlXDWI1a9FB4Q53pemDfj1mr55
DeG/VIT31FJ4A8qeW3hcA6g5Lv0GUuXyaIA9iXASKJi5U1J0ZcQuGKuqL4K3jX20
iZOiJG76UkDTbnR+ZNbssPACEl1TASB6XKygLWWvr6f/H9v/v9z0y18HlqCmvU07
hbsg64+I/vXMYp0EHXAfbHF3LLM/v/+18ELyYWx2WWamu6enizkO+16W5tVkDYFK
bAVQHff5jwI3eZFI7W2LmMFk7xJXsBo92ZaUuYer5D+MYszv5vrzP9bkPD+r+f2Z
ikYApKGn8u38QeC7nPbjsu0UjGltMKjkoe0v3FlvOpIrYtRIMnca/xyqmExaCZJ7
Htjtzu62NdefyBE0096xDyWgiCjmgmUlj+v2v6sv4Nj1NP72xRTjzLuRvu7C6sY3
omUiMLGjldyKkzuO4QHlrdF77whFw3Ab4KTTHNFovDyQN7SQYiuvZthtdy+pZiDB
OC9qr7mJJCFfawSdkuEKquvQE2TsgwJjQYebQVG7s6kI6C4YKrwhHT0cvPpH1G5u
0KldUBOUjMk0Fx/TQwLMsQiAqFmLCIJBP/fyc+lfJwImjTXj38u2xJ0b8kiLXMgz
XfMgwkKFkCgqSSuMg2dwG9yxMWFuaQ56wUpoeiFQR8TcZuiusPfFXZg5S76/sUAZ
k0YkLpTqYJYVVePGoMI6t8+CpDQ2G6oa9bWEuDW/p/O/zdBp+sukpCYADdE45HTR
k8UYZ/7w7D9h8xOOkhZuvqo25QSde3uriMnFekmKtW1DoZFsraxmDtIy89z4/00M
BVC8xiQfljrveqqAtoiy9W6SvKiCiwTM5A4D/MV1Ji/Q52WpZMGkkh5zlMZbvCGZ
eRR/IKysLGLUfHjjAJ8F+e3tlVH1E+iYsmulfa3iAkO2QuHAuidRF3ESpOD2NoMo
UnCYo1zYuv92mDPGJPbyOmbk1Zyjg4B7ZzU5FMHd7IVrykjmHRJTa2wEAe+DyQi/
RTWlrjwfvn5LlmkppjIB8wvkmrXF3reMPp+BnP5rdZUC6UDTO5wQYEax7ZAGwoFa
yJHiJBw3WOHLDQt8JdJ+BxUE4P/zFlbSsGxQ/cjflqdduhQbdu0w9gNht8oZO2Mw
h8GABWHh7b/tjxfNQVPAop5m2XfAx3imu1OqceFuga8Fn3CSaQ7AJS4IaLXcJnTb
qzF5Dr/PdlZw7QIwo6d1jrfq1x2hQ8LCWw8/FQ2MDodcRkccrhliFaGH4ajIxXR9
RogSZ44QQEin5/DOZPIzwotMCxQn+RcUopCu2ooo5BMKAuBAaoteVn3+pvICIwJQ
PV4LvggoANDHNmDuaQXUa7oRZNgLd8bDiickdxu1yF09JX3IehTPhSXjUH/bo4om
JXQQY2gy+0mV77zmtb/CGg==
`pragma protect end_protected
