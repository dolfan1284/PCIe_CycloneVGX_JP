// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:01 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GDIZaaCKs44+R5DqBRz3QIrmVuDvk9lkVhUIQHYOOrIrmmew1ISi39FwvcVECwNJ
qYyCZpK0JJd0/dYcAImHxYvhxe+MctdBJul0zov34PepjNwyI7b4Ml2lalEMS6os
pqJlRZwWe/MjK4YPdYlTwpapPBl36XmhfakoIyLmRYk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25648)
/xj3oy/ZsdrUiDFMeBgTl1O+SIRTyM07EBZ9NOPBCxsl3qzB5h5v+iLK6NTKRgqx
OVNpJxhJ3s74p3Ibo6agdvwR0uA82HDeh48lthSPs/+0Qy3hbR2j9RTgzyj0WLxq
iVFKVf4RZs6+yx9yRJ6V0YWWWZCn7KsY2KAuP04UXczwvnvHaHHm/2DPSVL5qdBh
SLtrB9n9s/zcoteDIDd6yRehBRhNBc6uKBfMwy0/EFVUeSPZ19/xsOapQKUhKYsj
9Wc9bmWN4QIj4f3nF4Ej0tobV+rKS2Mjci44oyN+c0+TZH3GbeTc+GbBNZXuxUzq
6R5z0KJfJ1nXznTShwcZ6LI8ik+m8eWShk1kmdyBX6KUZHL9oSC0jh51lQtRSFO9
MHnmKid2mer7C8M9UIGdIx2Tp0M60J+f4EM4jiWcbOZdV8vbXx+1mNtQ9NJoF513
vAMewkwsqB7fdC0zgMl9nmXi8RfCssb5wzq2YhIjv2rPuTG1HElUI4TJ4vGJ4zZr
6an244HuGLln23OFNRKlr/1HNeZhOgbEvdA07FcbxiaHh66fLUV5eB4XdXVMsCPa
X7IiUmprz6jCQfJuFvFyvyudgK5zQ9YkeCIEeQZ0nwY4qTaA0pACg24UwrCBUa2M
7rDdaR1rQ5agcABGTngLRG/gYIC3BXYz47NYqNk0dp+NeNDJexkR7QQE1Db9OXHk
aQ3gZD/YzZgisAMcE58V2ovo0TSw2flkUlTS0Hz5fheUIE1FgCdXd4cNFAXZLnsd
8JofeSvbIWXcOKRF7jIazk9ThpByNi99e1HrIE0aHVxFYjJyy79FcAv5r1/1PzlY
CxFFEcpA3aJlQeNlJmLsPUVEcok2n/MrKCPy8pDYNAIeKyXjTCvSXZqGQ2ZzJnE6
c3f3OdPQOPzf5ez9qOK+myLUzP9tPPbU2hUldmBlYua1Vj9FzUsojP6BjTJ4ZqLI
KEcH9KUX/InpfQhXk2EkVGuIO66OK8L2wGFAuZ5u7yBj4R67xS66SBOKealgrI5J
e3ogVKzCfqglG5UqNoUMrSxXfSBC0PqefgiE/++5RZgzM1qFAsbjcLDVL0fgTD03
LAyvyaR0Dgnq137GTwQVONGE96XpA/KNTM2LHZvoRup0Zy/+oxoIR6o5yUHkO3ik
ZYa6QTi8Nzmh34kcJG3/MTSriuPJ9EW+C3d1bMZIQhXI2MV2EoPeUJGfFjB+deYT
2rig9EbJ/piq2Ei/j3wiK/egvKZ5xfKBfchyIEBG484KancwDu7InHTOaU2cv9Px
5o8qVetAiLC++DnAVzOO0TQfuRrYe0svs0SbbQHbudb45r/AoD5NdDfeZWkm7AO6
145bhRDGlY/ZqPzaPgGe90vE7U+Rmj/UY1Ju0Ox2SaQlvJsCiyTBKYGPXjhA6E4X
5Ksewa0bHdF9Z5iddSyJOYBRbPKqy81MPLmJfytT+1F1SuoWGxnAKj8s0wStPbG5
uOtSqQVcVSbPhEoxjvs/+AHTMcml0LVWOrk4bcOQR/WrEFzlFJDuzkYqqjd1WQqr
6wxn5OCmWuouqoSr51d7IcU1OuQ1FNOMO2cv5iVwdLiPCUvphdy6cuUEmezEi7aY
06FGgCwor5TTtfXyDTgi1v4RofJ841WbPtnrJRSJhGwU88BSHjSiw0yorJI34Gxg
pDFkqajtpIXtAIWLkMJqRYuLDm0sfjkiof0DTrzbvMb+XDvE2QQzjHBYIFi4KFbn
bX79FaltZd9MaWSlVH2ANGCSCl3Kie/az71NfMYkJc8cjM+KmLGvrqmyHPsMTdUk
99QoKR436BUFg1qsMiA6y13Wos9QM8qn+6DF2KUyCmQlz5/tcud4774SSjROGUkb
vZ1uHY+Q6LPUAeXp9LGF2ISQrr5yiXhniYQmhfLgFswRwqEW5F8EMiZOeubXCIXT
rurQoohZ4aMGrdLGLF9BeHI+TnWAQHvIsWOgePac9zyXxpFF6UTPofZfjJKLHHXs
RLfqG5RLXn60GJ57ySj/32dbt0A4RKPk9Q7dbcgrx0yxZyhMHNQVRbawlAaVE1V1
i3rt8L1w7K/ppX1ro7pcxljStt7Ou+Y9CcXsGbRgKI7/cPsLUsCyrNPQSzKGyi7d
lMIDnJQxTrxjuzzu+KVxZYDL7xTqIt/WOQAQhq73YZkCG+20iUbneajl2TEJZE/k
4+a44hfbK3THGjU1A+TStu81PRgQ8mTLbayFBuU/7i/XmbMtFCMkBxtdgJkSqS/k
lDwdLhhc01BAsCdqxn5LgQBa1weEIZEXdDQywJe+m2Po6LZa/cRvOkXwVbbPb8tj
3lW7ZntiojwcW1+GKabkjFfIg0QSrqwzpj373u4fcMaflSaqwRu8WxksvOvrhUtY
Jui4bIV/EDPVABj532+xm2SsTnakXtXgdOgUJZHeJ8g1k3f0yx6lN9U6KWwaV8Th
feHzHul8Jpnv01byiHYREq2rihW+J+2D5lyIp8JJuTUwlKneOWWmOxm7HqKbjT8j
An+scPuYQR+tGQ0GNuuT3X4jIyqFX097Xdwje+X4Ur51lRZg8tXB2tFYMzWf3B+f
L03iBB+Z+stXI2rc64NnJcRkOD2j7kwHg/gHabYrTq0iNhZYUP5tPtD8BkkwBuSH
eqBmihuN0Zo0PcgH8r73ogD/ThiHu+AaTN/ZsSwnO1t7+4mau7Gu40vKWNnrOSND
lBkaZFutd7E1M8Hb6Wuq/VrN/0HHWcORqNI/AcPpbQ/HRmtBG2OJcetOZW9JELVo
eYiSB3n784ePOzV3xVKaWbQlNDhu2aQjK5zJ0wgHip30nXC6jGsncEPVHh1U86Ft
ZYHIO5aRKgh7Hz4yEyvNaNBNmC61+I+JDSuPPo2e3YdOzjtnIhBWDbw6VLn8Kubt
OAcr47IHCP/7Dmx+JOdS17qXwymhhvShVFCOe5VEKl4fvvw+FT3GmUc/jV6kjpWf
h0RmhaFnQ8t1R/ms8VkiQZZeUpm86XVnkznI+2PoXTQUlphrRo0LtdzWjfAHtxh2
4quFK3cSh+ZoshNqwPaJlXHK4mG8zXkGhWtnj2iQqFb2jkQWDYpyo39kX4gFvmGe
eAfCeIK09ISF9Qb/UxO3zQgXNlnDGBSD2UKd4ZwdW0eQ2NM6dkVcseR5Et41RI7G
qSns6Rg0iC5jWIkp78ihppQYnLv+5kwaeoFI9f+VZVpLxtWg8Anos7h56t8GYyaz
4OkrUStWcQMma/1fUNVOSx3ZHp8bi0NS6wM2ZerrR0raXR5t6m1nFuzKmwIgRmIQ
wRZ0o1sLAV10EdFCaw6YYKIWJL57LmPM3Dl1fdc6lAakWHNsD7Zc7rTsyU0HaAmo
DLWMTiY/EfX+wwpK0njzHViiGYrvIvSfmUHWL5Fek6CKaGumH28hWjIwLzTnw6wu
QBMMIao63GhGqslg7xwh7hIde5Ulo7qNuUQNx2O4eQNnBrDNiDFPzRaXLu5rTmkj
DZSBo/argL2l6ACU6KtLqWwKBpWG9PCVO9jBOc6udLvG2g01bJIFVAx3jT53fNOd
L+HxApq7ahAu1+FiDnLA4tEx0FOOzfAUpD5LHBlz0qiUbPXF899qLHs4AqOv/MX6
YJvJcNxmakcwx8gyaL/54D7HS/UtrYzGS7ytvpmWIS0YxvQ16ewnBWQA8J5K+jFi
t3/5GkZUwJ5+FoD27MK3znP9uTM3fP4TAHlnD9a6RHDxCdKBbUVx4Ea2KXVbTPE+
DUZGgy53PPxIaAX3YTfH/P+MmYwCXYH/owZK8r1n4BXGB+GYUH8PQIbmUwBhrvcX
jZBuNU5rNduXtwZhaCpOS5Yyu8invzjh0mvybJG1Y7aKY7efrPPVpf+8d6B81660
EA95iFi37GEN50BHXBUHjFtfwowhLoawU5TvI/ngJeOnQ9oTv1hLOmHg/lPItDMI
PODAjOm0H7a9hmJeoWLxFoVU7oVUUi/La9DnwOV/J5lzLQQNkBm9d5/ZmWRJz4BV
K7Xkq3k5ATMSark3jVvNGMJsMHcFyVrlEDERfZk0cheaALyp6f0UKJ+frNPAGVbQ
O3r70EjKozMZJTkBkZlRejmU+e7szdqFjvVbZjG3okDOakY827uoVSVIxN4+TQi1
IeLs6sPuCfb4mIF3jFC3M7QinEw3YhpYMG3v5fe33eHnAXxx6z0pB4NT+7ICM4A0
N/3RcxqHpderkhYVGP9XOIbzylDX+EiDf+lESaTr8ekpQtuDXNP5XFaRlPTgPscW
ZqrkNKRZPOIS/9B0OxhnM+PuDnRRFmYzAf/we7L+xHONn6bWJaQpfUyfQThdBzop
sR0K+R672dzADxuV3ny94usAi/Oy1/9/jFqAG4kabBT98sHqitLFwiW+IFR2nSDA
rjLmApGf6qEucA+vW1CeA2/pOoamIgA+OOBcOZHeklqGw8grFJOlAu5fAcbfEM/X
u+ejWkqmxpThefohyWnlUlT42z2dI6fsOEhhVLnCAU9MWgsXUYZxGCEmtHMNLt9Y
iSl/+3p15bI2EDe0O3nIhlkwM6TIKIXdy9XaSlMHOIi0Nn4u3l8L36o2qEYaQOaJ
9fNIeY81AB2XDOisswYCue5L9GGtKyq3cnlR5qqCPrJhVnR2dDc0MpmzMmhqARZx
y35Jwmp6Kqm8mQftH4hzP1p6aIxOE6+xEi3cD5P5HneY5I/J3uCLqs6Ke6FTnoLi
hKxsUN95ydYddCrAPJkILUQ8FrIZ0KOiF3vBAXvlIKb7m1950m9XNchIOkUKbibz
++iJ5WXWSfw0I1p5gSgC+Tns80Ws45wNlNYL/15mQUHwp4rZUV23MJF4AlXDDMsK
RJbhn7GiwyYCxxxlrz1UGpBftNpyNkcVglvc0Fq7cG+kJfvQCX1qfCERaLJxAKk4
RbRhrrv5Ux7xsgr+SOQtnJJ3Vay+XXt8B2XHzGRgNE9u2XHNUZi3YRNvKyNqdKMz
u2ul0i4Q7EWquzVPnPsLMN5nzcICthGWua+isELN8j7EjU422cFtQ1zsKEsOD4qZ
763ryga8AmTtr5TEHbcY5Rjh+g3WE92HYtg9mR4o+ZiGIErlGpZY0E0BPbho7b1S
+rt0vkBk0TvrxpvUYfs/cZOSd8SX8mXF4qP3BCFhDWk8DVH+X2LYCva3hkGVt+d3
Ce2v/C/XA3mgibiULnHtY7q492AkBYdmLcyxwG7zovUZtKlStopOeqbHgzBVfFjK
Hxq++k5jwKoKDLcTiBC4mGj1qraaUuOdPjNoYZXO+KzxN9VmpdxuIIxXMJ0aBwWw
r08eX188XSm1Mg2i2zdUEgw5W6HqaAFbyqwQ7UzS8IpbT0E9zGVv7ACh3WF3dydb
EpI66UD6iWlvH3YhRacV4WWkDuku+Z/hntV003xV4NOdXInYZvYxbCXPQbeUlGeI
uG2wcmJDXno8YR7bqcGV/dN6QVwWGRagnrpJFB48GgkhlBtaJUSVf4FhXZd1rVXC
VDqi7AlvRh5kalhiFTqHlQMJz8Yg//2hxNjZ32feX0nc3YjZO8fI3EpLs1fnIIEI
coY+XQRXNvcXmt8ih5eLR4cKAHYW6fn11jqvup5I0O6lhHfPuw3uFyHhOX37ARQA
hA21VV9Ts3MLpjtt778ScKHAEBAlzvDRsj0POurqSU8Uekpz7ca6e7tVA856XlhY
ShyJ9RQekm9T2a0izDnriQ+qP6Ou11rxjK72QrjpDLf5BBta2/zTTFGvG5ibwQJg
lNko/QrD03V2AZ2ZFRAFqjG95Gt8fZ4PHXRGENVbSeLKf8X/CwR4iOaqvsL4qQL1
aTUvqajVFKbZ8rVqxRelC+mX4rqJ3SySKdf+5gXiHxfccKmCtOoYzeI96bUxUlI6
R2ewITPmt2E/5CSXSTkYfySRMBy9jq2c3+Z1QBKru4+g2D+w2oPFH3DuFen23Xdu
PLt90BzGPXV4Etw67nYOGfYDpXa5d1zgl9xxaLwo2fMOGTFoleA8XaKQ39PALCcf
i8lXhCYGtklI+Z0fRbVa5ZXiSFRmuej7EDLTaEIsUN+jGZ17dSsH0Vc37BCQ7im0
/m+G5G2qvdNpi8rvXLiDxXgoD256Fjk0zB2DjSY879eQw+aa4vLFF/JTm+UpuQA1
gzysRUUWFenSpiQpW8sWmxKQH/5D1Bun/JWEO70AhfDQrpVklhxjK3klMenmxtKu
qf3HVohvPCMqUlLm5QlMuEtb5VrsmLp4Xyaly/9t+oY39D5Jh9audrqbwrDqa2k+
5BgQntduULjqBoBQowbYe8cNzL8PNW7Wi9dGY1ck3eJxRrNy9E+6Im+WNcrA/jZD
jIf6g8je84jWBBvaO9QQNMNqMd1fDv9Y8mwingEMfKV+DtmxLYJkW4IoT3C21erM
bmYWdTqP2e43jsgWFEyVIHV2AkxmZt8h7YvK8N0lUhMd9yBMzNuQB+kjbpFHwQMF
USzOPseDCBuDwPlvafqRBHWNELKALH7rZxER/p5Ije1pZQ+9N8M4JhMUmxu7HyFq
UbkZLcBA8rjTQkAUe5X8mwjyUPncRq9M+SL6MYPpTeboTsnmnh2EOpHPEYyD6/9S
1wRN4uGhEWS401merDx/bD0QMVbHOSutKFXgOKcYX/ZRdy2uR+nGbvX1C6mVIEKS
u9Z7U3Tu67GKusi74itSKp1xRLtoaTFMJHqfS4hRMLSh8SyD0WhUvFtuGDqg6wM+
KyqGhw4UqYwbL4bWRkt4I/FgmmclVNkg5K9ZitmKo++Ayl2/28e5a3T3w8CH381A
3Hv5GSRc+7YQ6EyWlOjSk51uGbEmjZnzd8OYrTR5jfsrL8oLZ0RGPKRkA4A4KbXz
F6j0lXTsEOMhNsF9+wotETv11TaKrpH/coxoOEysQaPvBkMPkHYkFEe+fL2GM9T0
pAWpo8ViYOoKLoRwZ3jasNf1PZCVeZvvJeQThwAq7GsjV4F3LXXKswb3OvKLgMG+
JIN4foR8+m2VH4NA1dHS6EQ0Bq0F0TmSo5RCGRj+um17dhtfkiEvA9dAoWTzVv7i
oU7nFet762RviPeOJuUHNBM2KQUAb31P2TCvY3qF6a6FhwJ4Nq+yPc6F4zpXdtS7
vvrA9eYwcRvETzw7WVKbHs0hm91rJclHTsMynWkzI/El0d/tgh9BBJE4Wo6Uqpt3
USJBkFtZ1xBNLnyMr3qN4WWwvS/5WM/n3WRemjzbfzPPNuGMAJjtlLmuGv5cpuC6
c+OauzVrRE8YEl/Gn1qJ6+9cH8sq1hiSpqdxQTjdE1brpLYjrGkA7GvvxQ42RL9k
9P2Tlr/VTW9F8Cl5Xni06ELEOlI+iIjPW6ggc5TuTvOmyCipfUv4nl1tToy8DgL6
fhZzzFPWmoVTr1L5SX4y9VmctiYAjovMV24uwaJ9sIPRII628oK1dy/L+0qD6NIO
HXgoTQdkROMCQwJL0DAxwXtc+RMBZbLvyrIew6uiyzTlClZE2d2iJxpn/L0cdOEd
NoWYU+bVhZx5IHt5R+Wq9Ss4hYYINBn0TYa/jT31BbhhL0r4ZyjR5+/IWJVjiT8I
1ifupAtehb8mf3STk9f4CIqzqvQDhiIOSGvROnik2ZazevxH4k1p1dR5I4IlGEvS
QFttLpXx7NrMilxHIci6wPjX1B0y7pL0vov6eoDyHpRq4EcKNYb+nE5JRiq4PFm4
Ar4571p8Tlx85jfZaIG2PCc/eCBPDiKrizntjJYny+SBfd1UpKuz26PkI2RA14jo
cnAVvrZIrxzIAByK6qrlTUIleUaCpEcPZ+4gBpN1QobMsc1puBy4iK7xrT3uORem
xuCJnuF/vI/vNi/ggZngkNvAIBOB9o8Kt77Eje3BrqWL3maj4XisQGkscrRc36TT
B5a9gp00BwP/VnEk399+hTT7vVTuhEFnM+0E3ORmjg8Ry4cW4aNFHEeXJyb4lTCE
56f9KV+UuasQSIB9dAMFUdeML3wSaWHcaL3v+whI6apsxvAZeeyZOSwLwQeNEE8D
ZDPdwuxsGEGtfH/mPchjOBERyrSd9HDIHG6mP5tAmJ3+JHLGUd4eDlHgJ8Ul4oMZ
U7sQsP9aWUtitCjqrBIGwsiTho7MY4jpbzdPVLAwhfN3b6R5vzheMYnz3hQ4cpqw
juklq1S4ItDAD2E+adGMcvxK/33tLJpbS9OnnMcC2n/+SUtPz5B9S7Ne73DgA4LG
oyzHbR8RDjiBRoM+kREM/3kjtlKu0ntr6j1H1XSVFRlS4mdTwxQrovRF9P99LqQc
9e8WcSpGydvLuW5/A683jOAePFAnnabYDWS6Sg0YT8f2SD4v7Enf5jmR2anN08PP
fOVOOkUmbMOEi1QZmd8DdmgcSoikhJyFRBmha8gR/6AT3F1Jo1TupNQrk+uhHAjn
XPYfRsiILyptKYl7Tj5RbM1sj8FnUnJrCn1+QC0jt1YVsl3izbZvzQhMTOTuJQWe
xCLyupp7f1BTAGftgPcfcRyMUyU/7dq3McPHDWmeR79oOaAItmplBOeuP1GmrLjM
RhL2ngZPym9TOIqyyNOAM+g3Xm8wz2xs4DzykbUsuOgJd7wuzTbz8Dzd3cxzYBCV
J39XMgsPDLA97fOvlyphCXpNVKbTjrOY7cCx4VtoXyUqIHV6YezOtRyzwv36x2Lu
rwQfuQQxtsRu9GlN9x2ue+0DgRAi5hYtYjQu/PehP4urbiQaI1cwM58hUQjQyabJ
cysDpNuuRJCVmsqeF/bH1rWXAKalLuCDot/SFhiKhkT5cwjW1LlziB1A0/9B8SvC
5xJFs9toxND80Qh+QO7W/3RXQrVvBlTBzir9BxCXlyu1QGmCLwPq+hXajjwJ2S4y
lBf7sr4iCP9hF56XjtawkTNhf5nkqGO7SoKoOX0i7kZPXNNq6qAp+uSOyTEifvVX
oIarKPHMMyxG57tczGJc4go/JKgWLSjGgf8OuCUJLUzXcePwhg1rKqZEZYRLxYFQ
1qK01bkWDbYJzPgIhDvwNChBPG6H13Re57lUezEIPI0oMV7c3HFJCHPnW4bweEXh
r3u7/SdEDTzaL63gbS6aPbuGEPx7MBkbIGU8cpWHpoSX732XeqbV8miT8z7GkKoh
GDvi8f3EqGVj7EwOwmeZ0ddIuqipgbqjDbd/KtY1BKSsIhbMgEpRQZZxggArFmhC
kXifTKsIU76pi/VgmjbMrMduFR8TsaoCDannXuopXKbmyX8OKCxbyXtCy5sMINet
jzQ0zPUn5BANl1fjpDcaTz/KtGd3SV5tkoVZuL8iQs8aa80HLA0GgW4MD/pplej5
71z9lreuZOCwulO7dBfWK5BeHZOOU03ZoUtlvrEa+5ly9gJXafAabXQky7yesE60
QJWEILpgWTv8ojk5hmgGXkPDCzFAzd3ycXPujglvZvFExYi6gKY3tkLuWUobR81V
o0Ejn5A1ZrSHVpfYyH8U4JrimpfEPtgD58/4/DRR5DGenF2XUqcBpRT130uSi7C9
QgTtoVNwuB8ZAWbG9SwkarUf59TdxYABE53h1HeWFVTO0CrP50FiDm/rcsPKZ8WA
EsTloqz2id5BSn3zCAfbhYSn6odxq+0RtVbHRCiFNmIgixcWiSt1QALjNX41PZzm
x3Jx7cKLDMmTHPrfQ2+1goru4bSPtdK4OegR6HF7rZYeInAFSeIbJBRQEkhHSUt8
5KrexOYD+fzzwYYxDt9C7LLmvVudrC6uOQnTiaEFlLKrHoTP7e5JHkdrfOFyo5HT
DpYWt/j2Z1NQi8LuoCoHfZqCVZqzt1NVdYOrt9L88sTL9Eo33seXSRm14aWhPnCJ
RHSsQ3MSGTua+3Ns4lWbeIDUGWZtKlLXnQ1mtmkl6UiwRxd3gCMfUxGJCYj0DDXX
ji1QTkXziOPN+Ka14UvCs5yTD1u1jmr5Cw+T2qLnfifVrphO/SFnYK6TP2SxsXNX
UVG97h9mllNr+PygtvFy7UI1EHRYmf5KjN4G4suW/9YVBzpsEUxe/uR7c7ZL5SSQ
u46qDSd6bqLMaOaSIy08Grl8YzQme2BujD6LPG7LCivMHA8SnhvDMZVxXFRYEt88
TsEsN84xY5xcY6x+aPeaM1a3reIBKO8+Vh4AL3xNADE9P8hwxbQMyNt1CRjozinN
WqWuwvoIg9FVD2VREH7GLH04YSK4cmQb5UFDFdjKGL82DdtaAJ06yWUrmeoGPBY5
rbfRL4JIkevhtMoh1+oxIqkK2Qb4aT4gKwWUtmhLkap6TheKHGbd8VHLN2+6VRm8
jhbWqEHXjUUu9XG1TvRXZCOjZUFINOXnhza90SCfbbjMYWH5r4NBX0CDSq9hy5Pv
6ACXFX/h1FQANlmZyoXdwhBIkohUAVaRVhjoprhGI5Hcg58DIMz6148B49fT1J/5
XNPFHUyeaUQI8zPZI0Sj/T+6N4pudkhTLXDuJ3jflxd8kUb9Kni0c5CuhqnkwePP
jRn70QMSZ3S0VmrczTqDgWBeDCdlHe5nCfiwYlTpb9elepj4wQc/bzZgFjPRcC5n
ojdCsGW3pJU9uAD85LuIAywxVkSa4kRWAdPNilhDQj8MsVGwBvoYeWOwcRRvOHP5
SgI15+eE6I9r9IHRIdAYLU5KzDRtO1gcKbyd/a/24oJHGi0wSt6M8aDhF5mTUIrB
5YYH/fthIrz64ONU7fjJiHMgWTksBl3vC0LmuA3NZ5eYYoR/4eLHoOLE2GWDsoEG
mmypnHyt+RDK3bB+RYH0FZX3vfNROBq7d1fELBEGDA90sHp6dVRwiXdWkprLpxOE
FIoKzdvTGFLjpyh7AoRrZLT8MYcS9nUwwOv+dgNAF9MhBt6WMGQCd5yby1Dcc6Sl
lHbYX2VcuMIt+R637g8jgkMflEKVX87Cr2M5ICz31EKhfWYH22mgicnHWcjHhiWC
D2CTBVAoUN+Xt5eFoJ07PXONUYeoFwF57mNADuB4JtRKl/BtJlH+2fC8sJX940xJ
gHdGPC0u5xWBVhrNPvXcWwfuQkBZLPUClhkc62uLOt315PpQaHHJXWs34Y0IIEi0
U6SBzUXhpk6ViuwO2/iDFwgWE1N3R0YXAB8z3vzYhaiQtM0yfxDVOH5j0Ab8OSoW
9SU1taaBVGWWDWzJlEsRWVI+5YgWTfCNg5PiRDhPwhEncTq7GkVfgcGQsnNoQPOP
nkQ0BMKSbLULwyiAKFhvweVRXjiDofGQKH6qknEQF+SAaOJavaYIVINThEyBbyIW
pTQkV+JEPivPe+aum+PaaYV8QTTq+j1IP9wXz4DesXFFZlz+A/eKPoohD7v/W+bc
w2jfQyWk+cAL0KMiQ5boY7aB9ow+mEs+7SlNkP6md/NLdQSO04RrecuV2+EMnTiO
tDEkHOyg+kH0M2dcsPcNgd1pwk9tIswzB+P1b7MmLLxgbm2h9vp3C9Hewu2vslRJ
ZyrrZtmJ6gQjLuZabfzn0t/+u+7vBRDfwGxjm3iADYszpNNeeN63pqoJPTdZ1eVH
8uYBiYB1riaoy6CI50/F6Je+f6tk9B5xWNBnqbPUnogIzLhYnlcEriMT8oyWWO2X
hwauesJEd/tuHPfv4BcwcXUo/lDb2qMtgtWqBIjUvIu1EOk/AknOIoVN7yv8zncG
qjl3CSsDaENcLFrNVLNoWI/Z3cg5pH8q8/rynJHh19LGCuwHLEm0QeJg8YwlLCj3
WzmqsaqN6mwXO5DGVU2DzRdU1JHuRjR127EKJSgTxLQLm1zaeYZCZB8UACwCOhu0
nAoQ6ediNmmYQJtqAqdAiNvkTrZPhfcYYlQwB1IXwnLzyyI/1nKeT1CKjJqeJ4Jk
k4B9RbaHLhH+LwBNdAL9wgyBhHw5kSkd+QXC9MtleyjUKO4lkyBOBfuSfzs1vvVy
KG/G3aY3qmi0iTZk+R3VUb87nOk6IWRNq8KxggnksYEkMf4NOtrEL6hSn1ks4H+V
TIgRj9CXVKmTVHwVV1njJp4WM2jNW1TmPOvaEdUnZtvpOdYwpILAtOn37ZzBA8n1
PdU5U5QEpV7HUHmo5j6qBPEaigiHM3ZKiK83EMXYQUpiIj/sEU1OemIGFnqL4idC
RR9SJzbFcN54XBcg/2bzFeeCyYv67VS/xkmV+Fcc0elJEUUgzlao9TZMhrCWpgPA
vk9alAb2XyGQNuDyepGmMidJs0JnxyEpG+qaJ8Xd7g6CCv2xqkIfIor4QMI7G21B
zCtA/4k35jdkYISVlYj99dy+YC2NDQIZMR2oa3f3KvcxvcVH+w88YEYCz4PJSAoo
ONyvZB60RwK07jHtt47iomvMme2x/mR2+lGuEbP0sFJE+m9MYk2QBPSdjE5qzrUf
zr+93u5zse2uFZ4o1x3vQ9+gbn22dGxpazWSzCMw6vjQgkkBpPGjoaqeV+SgypsC
bUy6YZ47MI3dEqioBIRiDOMgLamZEjqpM0+ntiEBPsuPyhSwD2/BXCzO7as+lmbY
emQkgjybO4x0XbUtOp6xfW+n6nD/G/B3d5D4GyVeC+A07x8GdDiRnxLsE2yizkJW
kY7b2AzJ97O3bu9PX7uW32D612+PiGlKlyVs2omiUKuE0NlUnAzOOpdM8nR/Am/o
pAYJGR9OaqE2OFNUGcQHNkgchAuB/SnDjONKo2FRS9BoU7pHvjkvvtAN+XEDh6CB
/wL+I/AXO/lN7sAVIPBoSRLEnFXD72S4epD6bdl7w+WJLHrxQRN2U3tlbeYzD0L2
1mlz/b3xvUHQTXFu3z8zu/ZtlqoivghNg5J1WT6A0O9XiaLD4WUuUyY8ZOkUiOXz
+hrVhPQ24MH6LcCxDnl1H3mzVXUvyoTyCGPOfAeEct2oLfrmqnC3qyY+6msMCed9
vobvKjvAHNTDIbB9PWp5yKb6sCCf6dHxa/g4xk125/7pugPCR4Mf68v6nrELi+Da
Q4XsSZJn8VYn0xQzEhJzkaitksMQ0Zi0W/3xWp98i2kwzsBxDwKP+IxmMOmGPdc4
+S9Xl0J7IOZAx/YA0CkFnxWtg4B3AxW600cvXb3+7f30/JeAKwq6qETsEXPpYynf
WWQe7/EKBx9Ftdgl5r6D6gxOUWne8mcyOw7VGGPJqGISCTAuEtZJ4qGpFK4Gpwth
V7F/swXVbhbDD2A64PD1/0pPGrmRg+WgoebedqI4mwxFU8IzjOuq86QMN4KWThaz
YGSKzb3GzHSGiEA6iha9Nf2rq12VzAsWXvI9k1yr+vYHR+XcQJv/SPAKqJdCTl7K
Xj9Ii/jc8DhO5Zrgh5L+Agiqq4rvIrMg6h3j58bhtDvUJRiktFQmHSxFOBpxj3vm
U4uposlIFy1fVjytRNNM0+mmrM1zRpLOUpH/E6dt0A08GtSHUS0Rq77qJNldp90o
hIKC5cv511/Kq0c8DwdezNMuOaD/QgVgsUCxSQoBDon5xOTYzONkLmOBTakhJ8Wg
pBNQNbH0Uj7M0eCWY2GmmFN9kIR0qusNvKU84G4M2Xay3WhJjidWmgEatj0dYrhr
O4K0N12PAm9hq/9/+CU0fWorai1u6C0yhC5HXksiHYQ1oxOBozWKIs9pfOfe0Mch
tpOz8eBiJlUkC7Rnx53AdIp075qojl9Jua9/ESJO6db3oBOSd/lCinOzYHPex0eJ
KGfdRr+ySuJ79HVLWxaApnCHCLX2jvemwvhWsGpz+BJq+NWplXvvAPpBfJpCDV5j
jMOVPojAYlgJD0e2LpOPyPm9yH8tEWTCwlhqVybzOXxrBvZQUUBVdPSWKxOsZLt/
EtWM5nK6GDlCFXl+Q/Cy5vdGMNfhALzguEfZmUWAXFTVKtlzLtyzSyhdoxc/x6LK
fMPjfd4p3TbE+jxI9LN0puJqLU3vF45EpDZ5SCxASPhYMCo5LzBldxOAYQMbaCMQ
gnyWoBEami650GZ459XRxxj3kJGnstSvizxsCIZp70igThcynRggUKQGVRfAJJnz
QxJzT55d4v5IEqWV11MI4EwX84X3CWiFTUlQRKtSEIglGdfKer0Jsdtt6rFXATOe
S1i9aTs63pHM+gYfo/FQ4rBUuaen0lqot2WxFhu39CYVuzJA/BaQS12HngaZwMOo
r0oGZ23Jazo4heKPi1G/kE0edRyyzly1g0nwQiKorlkIE14HybFKCUuiQcB6bu5O
aynjJV12QaxAf4NjLRpO4CCJjoxiKvBAz+i6yoxjGHlt1r5zqhsZ5wPwYwH5/ovF
zVIRWtNOBPIVBeVeNYOULAN2cu8Or7W9wFAcJSRymd2cl00+URpRz40s2xWMqU8P
0GoB3abWbNAaC2Ft2B5gRcXh4rNFJSqZNmO3Dq8NTv0+k1mS+LAMXlu7m4r3Jbx9
ynq4QuFfQSDuKusv0s0Xb1wLl6LG9WYp1r7bxt6AFK9mrHFcIJ5bSIHTsaKtnORU
r0Y1PoN2jFHjbezmVKtbReDvi4xhOuxR3XYzu6bEBAwsFp48M1IcPSSSvS2+kpiD
6RBvqPIkubVPWpLZYXtsfavOOHPgUxtnVVQ8dH+wIJ6FnSz6htSvFt+rOtaQTOUs
C0iZ0LHye/fO2AdxwFnrcVH87ACBOQNBukHWVvutKTHPgy10vn9NB59xOLM+EAtt
hJR43nwD+ZrjQZhJz2zGJOD1PqtK8vkntlaVoMkzi2EQ5Il+DM3cj7l3rklPldEJ
lRO6cZafShTz3ONB1Bv8KKZ7S9lAtTSwhEnYuC/hZtdxHvu6nCdXCMtbCMCy/cAJ
f5eL9RJ9TQ+8BfWIrt2n2C32dBwUDhkvE8IGDjkZau/HPAUxHbe5eRvUdlzPrF6a
1VZK9I6A+63AP3cbVY6LA+SxDTxOsa+/tnLjTanT3TPX/8frmNDpu2it6aofHtm4
c59dByl/WuWBWcXqDNRsZSOXSBJYaWNmNSDdUPMvz2Q+8/P1lLLEaVWU35/QCh4h
+bAnu+SNTzjacDUjf2R1sfgFr/a9YIXcKUNcChXpxiXgFCd87KnNJPQGxF3XijWW
ay1w7f38HnqVLC7EVg74QQsFBwPQVB6HM6FWjBsfMsaYBlT8EEBI9Fi2gcdizXay
rzKocysAzYYN7J27GPYNk6cwteIfTB/soYSkfeBVDEZRQU23dOPfPO9n6P4LaqKC
Mjifk45kJiOyGmy1XOrEWpmeFxWq90GG3JG+Q69FBxZRH6uEiLGo+Eo2glorrH61
OSOYDlpNS1T7bkyPK9RyugVo4ZEQy3cXyEtcYjis3fULDrEgCiZQZwFw1WSka7RN
gSk0RYh/bQ2fhKQcKNVN9G1h67mcRbJ097dLtA5n6hYDuEtNJPmnE07PMHlbZ1ll
Ux7sLWT23vwQ2OuxRyKS4yDxyp10mFdkPNHkQPBcwFoYNnvSUtjSZKHT2YYUyWiI
VI10zkDM7ovgpEFOKPXqOqZjL5vEQrm/gp4iTA+uBBoB0yIVuqiLgKkhdNEcC/UG
Z8oDtwW1o6fS+wdMDpEUucWaSsiLAkkDLCuDRvcNZQOOJAphbP9rjHuNcGK6sQDd
MoVUp3+Y/rFy4OHDkS1vxkcVcnmENe4iaf22dYruP9K3DAbIkDhGw0mX8d2lBC+F
EV1VcK0puDrfL9nzM/CeEb86r4AEVgRB3rqWWxV//D3+i+Fwutn77EY2gInYpsxA
MC9R+LFxX9ju7qr4y9HhYc34v8+sF6S8xo6h6OqGjMsXegf8ldt/vBo9OMbeOevP
Gk0Ld+RaK2nb/D4DCHx2XU3+RFHBtHfor4TbfBh3pHJkcNAO4HwW1frt/bnhM04Q
x3N4zAingq2M5IiIt7cERVKl5E6joLnaybig4DkcrYJCUaYZkZCRUZciloYETho/
A9tF6TOE6T7T1wc/VE4zc4Ya6U7N9zE1RDsEXZ1P2HOrf0OMQIyl3TeQd+fQgvAL
HZakm3UqCBReKVN7GcgAjjCQXAVZfovCMTNxYEtAgK97frxUPQrEn5a6gkB7BYTV
8PBZpiwD1nCMsxZMRYLdlyjLU/RzGI9ZlheW+xWtpD0QjWl8v8NAyRzH6W0q06ra
ALk40Uke9cXPMeHjxuSHdJiNy7yZK2/Nsa90B406hw5jtazIyyFiyQ7QlQ5ipVLv
7fpAPVpBuOFEanM84GUAaOodjEt6PikwK1IfKmiJf+BVnmgY58QhU/lDuN3B2HNS
XOzG+jHLYT8fcgTeEosuihQffQo0fgwmJGkM6+ic4YQVnYnGZYaeR6iY3PPfcVW4
6xZYFKNC5UlhOMRG4p8vpGUw1ZWBeX/M9zktGj+kC4PmAHw1i6dO6CDM89QoxSDc
eO3PZD86E2Jduswe3pKhR11Gi0ML29HviicoanNbepIVEsjujylwsX1kePfcRRLM
/o8fDG5VtF6hAneRvaAFFi7opbMzpC5Kmn3Ri9QwZMSPRWUCBAV8WoC+qQB7QMLi
A6zq3iNoxApXsshMuqQl2/aUaVZz/KE5c0gwGr0YJU2hKhbRw2MWassx+wq91AW8
g26JnW1q1RSHG+kQXQrpXiiIBvB6fHPESjufWzOjRU6FrueTb7Ai2Kszu+9WRfjw
J8XvSpSbil2gcBMLTsUHeBeFFwLz7/I3351Sh6iB8PuJ97LBXN6GkSQ/eMx+k+tL
rklzcugwrlARzb8RWL5Zf65Gur2jA3AMSPWPaS+EMEDlJF6g4KIWjukLyjg1OMWg
b0Wsh7owRiEM2tRBXc2hmmN1C9GCfYmjYbwT+H4xuTASkVPFN0a1tRGeUiZg+1Lb
9fmimEv2VqYu+RXLTUDG2TxVHL1kf5tUdXued+OJ5ckNwJ2K1pRZpLmYyTmeifSX
B9yjUpCTqHUZVnwBM7R+Cp8VGPVDRMKpFUEBGxUqe8dR+eKzFDIi21AO5eROOgX3
K2Gjou6KdKgMznAvb19eDCSIVWecE+sfYXB2CyxNdrudN4Y9AvqgaqPMgpex4DV1
AsATBpwsDtr1INWn4m2uT91PnPQ4XXjyFVL1lfvzTEmqUCHZItcGEf1yKbvCVcWS
tsLcK5sgG/+r8GY+HD9GI/Hoc2hRSQP9IKYzUy5STQr7MqnHG0pT7XbeEplAbNKo
JWBpQcSSaiKOUQWowpPG1vcE52CPQZMJfGtcGnI/7xjC9u+SNE1CCe7lOr36GLWc
mi9bD8J7mPtZxbemuAc4j2VwmB+B/msr6JRdcPNnj3oZ37pFPb+3XHS3adFBDL1S
DUhhvQ9C/FyYR/S7UThOcPgRkGnqoiOfmUAjVsoZemEdxUalyQVKa1DTVvjQhAdK
RdHX5ueC5tLMzfyd5O5iF5FgtVWR0K/2yuuGgOBeXNTc0jooDns+AF70g5h+betn
0I8yaYGdmFDYDUGCtGPIxvQJMTWA2SiTSDct9YZFl98fXMO8Hkaw1gd63D4V9OJy
9JZokuTa2VfPZ9cgIWfsaTszHO6dkz+sCrpVnQ3+1JCZSeHydrMHMbmjN+ngut8u
2gXp2upj9n2za6T8ZbeNr4gdEos30sHiiWarbJlj455kg3CFIXp24IP6Wt4NHQxT
JkQgusqHGtJzDuIYawcjL4/7+0PMbD0tiS8xQX5Zf2XOOgpMWjxujJ4rftfrfW+0
1kuejT5hbhepyzYfSV2FgW6z72sysnb91qv6JBMljaeD37+dTIyoiJEEfMUXhQwL
iImZYo6Fm+wNMSR2CGPU2OHcPKXaV1F78e3NS9qVTrgaEpOuh352TitXwgyXkaEi
jzrg0sYI+QKXBAICtNhtm0kwQaHFF11kxxD7Ggxc6VEXSBRtRGueQOnM4AZFpmcL
TUqjbpdFSh6eRaprlzWH9oyyyyqCOxUTOpOnSDkwUG1pW4DMwKfm8yHHv7pr58Fd
mJwJXN+Shd17NvdQrtY86NJv454f8IUOo9lpHFbMURX+CFOrfTf1uIt3e1inav0q
Wtb3J7TDsQGRvIcFMZ6nRnz6hdBEaupdcIEKJkOCMXkb0j9jn4OETzC7FvwcH9c9
nAR8/Ok1gsVR3mSmmy2LCcf87j3OtzYCXPBewTKam1EUSC0ZqGeZhdXV2lHgsxgm
JEwi+18eADhtrqu00fFqc3qTtix96YSijMvUAoG8C8wbqtn/hjf0lAdAgebUa5/e
4DhidfXOKpOeZxLsq4eVecCnqnhI4sGmxybi88F2NAnn3hhngRLEKDxxUL8vSDEN
uWq3+vTVKgsl5dWoHvVn7KFcO7zrw4dTXSKh0Z1Slv31pPQmByENwuUku6IjSmO+
7HRo33UHAIDfIxjlO/ZaYjRNcoskLKfgHtpHy/CRoYrS59yKk7TIhBWEARrdUbXN
kPiTRdUh8F0N3J8r2/ptbRw1UOQ6H7mSzTojHyE9ON2pNzKZkI6Rl1KDMQezzUhc
2Irl0ph0Ku/PiMWhxb6T0MPxY/nUat59icRLFhN2KzP/XcaVTmx9eVSWTVtbMGn3
KA1ymNvAN4kqRc31vpbaIsK+9dkzJsPmzeKejFyTJYmrxytCcqTQJeV5wgEMr4ZH
1oFkKvnTzs3u+d68LPaP4nU7NGtGK7C+7MrSwsgh+4mtkhAQcPTJMgYZ/f3KKI1G
6B3NpC8+2q1I8L+eyI4vWeOZKqORG16NoOpOSMn/UYgSa0uUo5Tvy5wetQgUfnKQ
4nlNDAYu6/sZya3etLbLSIhzgohB6jG4YP2micUST3hqQ3za2YEyqPGMXbKS5oQv
tW5S8kP0jL9QFBoH1UoF+L+RI6Yl+F6ZysJRv0UccSZSUdXBbQGB03T5B2LmLz9H
MrEyOsDVvZ9wyqBh99K5QZ2IqpGWY128t7SfH/AjMuHc+b8pHLwKFfKd/5k1DJF6
iDhIjK0cpxJ1DY3c78kxV0DZvzyguIOHDWnLmbIg+9jANkz2baLI/F9PSj070P0I
329du6GNDvmQo3atOy2Jh2n0HqzJmuJc/Co8gJQ5CJuX/f+4GemLE8KsyBYY9D89
nUp3nBacPx1bSjXQ/x70+UAVBkLzBxwoutLaPCSDdppWOzjGPqDepIyZ9J6oB4SO
F9+OQg22/MLQuDAWwGPqX8w9oCWayIOBfM50C5x4vH2SH5Q8GkOheF5ubh/o5+S+
xQ8oMci1g5LTqCx2dzSKrAz7D23+XcPD9Nz9IdwuNqI5XmsUqJMshZp/bF0FyUl2
sXXJMcs0oSTYsbHqzppM5bi2f+1ZvpfZy6NPZn8f6qyAz2c/x1j46nbAWHB8cVOh
oZ+SoSDXZwyNVFi+7FeNa+pUByznxuDV9pgWkB4WqkP9PT86q806zwhP4g2L0aMI
lsEcT0m6De/hnYz6ac6MCzGiE6sdrTG1vufdjqifnSx5C0zFk8I+12w+z/q9pqpK
g4IDkRULH/jukMB915jk8mgDDa+xqJe5JttXb8mKPuJHVQ5vc2bXMl8xV7hhDNSs
ZSYUjYclx3aphxVfio3VosRIXySbU6yrSFQ9u25vZn+cRgchF2VKcum+62QScYnE
8n+2p7JsTJrUTZD4/XseUkXcQMCknbRfgUkf0MLI/AtTe7P5Jj4pCCsqgHVLoyQc
4KeJ5OJ9nyxEjlRzele6/xm3AKRoJFyXUczm7F5kXozTmE4eVuHVxI0AT73NU/lX
j7oZTx/I3p+8fwEL3KZUYLhwVdoBqnkHIcNa0xY/VRKulcKrKzv4UToUMysT8kyc
o+4xU32gEZ7T69HCWuoxn0QruOSqgRVSIVsXd2Q5+t0InMGAH9aYbIXQzDC0+Zf+
byGcQsGjO4/UJ7NRZnsvB9sA3Hd6b90qHwfMHxMurSaDRg7qo3l7oMe0hDn/HYj1
ctztHHCU/T8gke8DV4h1NRRn9U3RI4ndlA4U5vPgCccqAUmvrGST8O6gxffmQcI7
KM1akkv8LjC3/CkE6T6639KNogfORDg5bLZWPayRyAZwtQQxKzlPh4yTxZUYJ4WR
WiL1USGGx86YENw5ELwGjCKbPbssIzIsT3AZ+u3ZoQ6zVZ8q5UmqZ2CHEi7y4DT1
EJDl9dh38cID4U2B4T/WwsYFDiSOIuprH4xrCC47JNA9lTBFuohEZE9cpCyeg3k7
6tl7l8u1ayPYEdo/SQ974V2yyoEswn4SOEUD/2UrVSpAOCeFAG0CbfRJ3hsIiyqW
D8YbapUJgEj2j2X82bwq1kVCqT6fUwDstkotGUXaxYE1JMEUkIxLSZjNdFkpzizc
YD6JQNB/FcaGPLX8oe1rrB9HklshwgN4oL8b0G3nWfz055xGo7oOT76F1PqJOsBf
yx1uNsuvwA7+ENrKw53P1G0RdChlqvWfhWWgu8pvSACnbGH9F3Fh4NN5fo64GIb5
KqKoKssz/3ALFJsH6budikJ2BUZwwllLW4HmnA55cWp3uReFO1kODLoaj5dDLTjl
J+s3eC0nSrsjXHsSLinsnegzQGf1NSzkyM3dqq+gM8158yP6Eyf/zNWdKxK6oO7G
fhdCPT/kg5hlYNeri4pcxDfGq8pEXX5yI5JJpLRM8xbdIGpIImImPaqMS/3EZ/94
A2zPE9szxSMGYZovhHOg10YdXzuD+IeSajWuNtl/Zhze05I1Zab0FlQ1e/TWVByU
qPLe01QgzmvdPFzVPHEhLe6SbQ3DNAYnR56lhjHeCwy2HN7K+rTdYQEhZPvKnpnM
30wXteAmZkK3/C5khMdHYOwKFBWatX2C2vkWxYoxA/5ZIdMdt941PB0YYNmBtRR9
4fSmxMrDNvmIwYafHKARUn1KfNh4wQmqwXB/lEy/Ym7k3c4CBzolKSm28CGFFY4W
ibtN86Fm+yp+15d3fECaBdGkpM4MaIYAXqiHReQdzOd7qO/NLYPqZbiD2HmGMSYr
/h/BxFqYnJ6cKy9XYF1IAq2qK1QBoN4zn2gAlI6HQLo//7zPa0OaNEHouPVv2xEV
6A3DJgmilple/jhvrZ8YVA2bdc8XL6AywBpBkNeA4u2hpg0azqpLdI97vmAdirok
JwSG2rda1RcIDyBLHNVNUB1SjKk0vp5kjHo6B6LQ7B4jNZPRDpZ63+Hw64lq2Y8y
u09BIly6g8cJ6f8cg+FXhti5vO0chGWI+lXJRmUmhC5PDjYpOBKNcpxzz3TMQMYS
rYhmd+3MESdj4AbAdwm2iUdHKX22Le1C8OPHhVU/TDpJ06Q6isCT+Tte5t1ExpZX
HfIHsyCEOxfR4m+WYV+edDgqfIgio4gK3FfZfwakV3DJi+4xX6wlt0WoHlsp+vCE
IYeACSfv5RNZmNt5be8mCxDXEDjGaBljRregkJNzV+EhZkWDJqp1guWnn0NITcyE
DnySRJptSlaMsxPlNNUKkxujrZb7KQAeMMrd6J+LAhbtWtMsdFf8WMOezY1CvfuL
49C/vqIKggS2ssn7aU7yuI8PWhttCgPihy/917bf/+L9OnDfh1UJs1qxxCxauGuY
qTLoIgq3ucr4SSAQEfW1+7HlFYInynFlQSm5rptbp2iwbpDgoJLuWrTb5F+9Yrbp
jTtciMBNwl6EYpFBjjZIOkFQ46/6osSOmMNR1soEYt47i95PxppWoV6PmVpRZq1o
1s6rCXqACiumB5GLd1Q9hULxrnJZ6v30CTbLgTOdFW4OeRzi+rRfNMoRdcNDG2qY
uScHgnxj35pjb1Ee50P63W48RHp+Z48DvspoGGsevHJKGk42VdtiNy6xqcbCE7ku
f63xm2183KttQ2o4HH3o1NBrLBHZc+POEsxVaUpCneotHrvlf2UTWQMI6REraqxC
K8L7zZJzmzcFe6A14KfKAeaotzsKnU5SURFz1CGnmcnRmCnH8+SYDBb+7CsrrdXU
29S/nr2G1vS77NK2crc30DgZAtl/yDHnzwlPDhhbPs33Uyn4TjhEklS+pz9HH9Gn
2v9YQNmfV38LVIVreB6RBX1Es0AynrMeG5DF5jx/RAKlVp++yK/Fx5YdcWRHpI67
AnxevjvDOO+bJ/9HZbPP9gHZUEkEtAPQMA35QYTnhpxY5u1JqFEgQRIUvprkUEnx
XIbbhfFS+r9jx3LoyZkaD5fxfDUF1wZO2R6zFq7ArlCLLtpeER/hOcKW4W3H/UHg
TB3FJoFWegnGncl7QnLfouppBsXr3e5Ewf4g/hOUHrgCwDtcU6iEuzXD77gSIrYs
o1pR2Og6Uvl13nM0W2jr8sCMByIQA+STtP2GuDiwktfhJboiwt/T5F06l4QgWydZ
K3vIazQYzxXlIGy+g1b2AtZXzn/Kuj1hR46kmzqdL2tXwqYssSkDYS/WrYgSZT1K
ZDL0hX+l4ukWF7kUwvZ5xv5gd7CIoqXx3Rymx9nnACaGtUPTDTc+C1AfvcSYe4qZ
co10ob8h7g6jldN4AqyHBLGKlZZ1CV4rQJW35OZme21qd8MRVCyVC5xl8/lKMWVa
TsT/2kNrkYyKR7MbwTL8kdgQ4ylt/pM1wDJ21daDgBT36krvg1jMvtNcc0xIqEk+
hrlNO2JTKkUPOwYvhUh7scpD+pJNlpdGmoc5KD9g2wxJU51StFtLVHFjbwdDB8ub
y8gz8nY09v1R5BYg9FK/8KlDg4ENjK1ukvjmTGHyQ5gJ59q+NAjPJbxCgAOxQjL8
wwggTsqGU8x4wC4OtqAs6N33kmDAuplHT/6T100M8K+YwjAJUxAPRGBBuVBckA0K
TUrMCnLcEx17u6mm3i4zaERLROGwRgweGAinNU6peOKzBK/J19pdyNtX3ReadhXk
ya74vOKtik3NiVBXH3wDEd6x51p+k43VCqmy/6Kf7Tdau2lIRx67wxnriElaPsCM
w1DIPnCmI6Ll9fXsJAJVEyRAtW1I3N2eTIUF62qQbaK1wfv70Ep4TqAPMHt1ti4H
ryAA9Y8c62zlz46tZ0LoVLFJUeZ9IIkT0wNTnU1w7JLoLUTgSlVVOVa6p598hIWx
Oow74HYogH4IDA41LiQbA4aWZcHRQDnATHAdEk0Z2/kWPGg5f8zoSBdvugqE77fu
XyCMbXrbAFxTiBufIZDDweYgCaXzloYmJ8yT/D7ukhKHjAAQlczNAaEiq7wQenZ9
6B7KuaCs81v0VV/GxvYHENlFEhbpSgm5fH2vsWq6IBRqFZvEZ3Q+6Es5MBwPle6y
rpF4arVFUSlP16voWqmfNKQLytX7nO/xuQX/JqGBBlUfs/dWDIHvzRqqsBSGlSc7
4MWmRk5r8dzFtcb7f3tFyZcxeGsgYUEUi0UvvuEp/p6mcrdZZaX/DgJYXVJ5x7tG
CMYJgnEnYJmsFhEkgJpyaNZAgTc6aT3ptUzwafKhiTXCxBmvgAEaVkCyvB9w8UgG
+yDFnRUvi6Pd1gI+pSN4jwsljP8yZIq7wRPIVFgLFJxPDcsmM7LSXv6820Ptc/Dl
6Gj+dNxXEg2vujSLKKvidx49kEx+m14Vn0BAkVd+m9/1xwLPlPc6lJev6j2yp5sv
bkbSX+vBEa9yHtMkzJLAO0fjZ2vvBnWmqkchL3bahS9z7sTp3WEcmupKIEstoQlR
8lr+N/vXmLQsM3L+Qc/jLUgnb064U6QXQlLaYjKCj26O02Z0Ztl1zWyj/KzbhylR
vhoLMSFQRsanwapMZznTHOA3amPoaV1fPjZM9+nWcUk4Sx3kATWLGmS0V60Spi3U
kzdCecVO4A18XSmp/riyBN9Clw8r2VVtrncjkr3mQW/v+Ifk11NwHvdYswgKxSnD
VP7KKd5zM1u2CU8yIheNzEZ5FHGhHryLT8yMwo/E9j63evpFYb4EnCnb61rlTHWM
6hC7IDRvz3jdy1GDjN3BxfcH+HnZ7ceS+1XqamWyFo70+75o/ugs46lTuvgF5qwg
79DFavL8EIAFiLx/E1dcdA0Oh2C/HfMn+dlJupS4VnnVq/naOfDQo4ZTJ/Tj6kp9
MBoz8Yqo0C9W06zvo6axiBfl2LRqgBqPs/4YaMvsEXeqFjgca28klY+ah+A0v5mO
Il9wpwo3K3yMo34/e4F7uTB+geUsD7ARj9a0iJ1cR2BgIdXyJE8bSvz1gBBvwwyS
VP0Y+IO1de9VI5Tnsm1gqfvU7IkNd7MA2+5MjpQC4u3zm+e4aG1Hr7RfzWyWcWMY
nCJzdNaWn8pXnU2Hg9ZlN8e/AKw0+mh1OeVOuNrf5ZliwDMx1CFBZ+R1M4z/qS9O
rHqWU5Y9cSyduaJ8KxFa5hQO5fNE3h7ZZxWHH8/963yHrxnYN/U04RQrv5RhZgP6
/m33UgqZXHwjV4+mGo54G2RCZzXfyJS4DOA9untlVElg3jSKL0FxHydDh3fHY8mJ
ULYx2KoFcuYqQ0Oe+vaPll/uDpCDnrBPbfU5ae3doQv05CSdl4tA0aQGMDJUYxJr
mWB11mnbVdOcz0CWKn4gkKxCyXcSi0khvGo7wrxSZd5PjjrCmb9J9DcTZMvL535b
P3PyVVoWh2GJbtdHg8AGDjDgByuIFe6HKGHmhDwE/ItEA3KG3hkfcwkqvDX60Wzu
KmuJnLSYRhoJvAYq0et6o42AUTaYOTNtWxfQuCOit1Sbh2Nox7Gys+QR6QH5nvnQ
kjfK7duSV+cBxqqEuZzf3upLMtufq8umuNJiZhjdJJSktEe4QiFjk1NessI044uV
+FjknYhcCPt4caxAEPoVm8Qxjg29rvKp4JRDlNqvSjpE5GViv/fcU7jiauv7QV3Z
FdVsWYmBg8LdlX9CL2IRdh6/7wVnBTsR/2LQFujncr/664HdGgGYp4d1QnYJ3I98
QnNiMJka3da8YQhfTyzt3k7uCbENHFwjz3tCFjWM6e2QwL4+iPz8stLtILTGUalg
E+Aug+GbdZKyrXC8RtRc6sDrO8OWmAvHsJdneWkwm2kJIn0pqkBauo+iX75SXpAx
lppVtAHb1iqWJtkKZK/9vaNNGWxn3qGyNWn0nFHW048whtRiFuwvH4Vk36QV1dQN
uO9TaUCgD4jUwhFNlvtqMIyAo4M2jydhJTTRZHNWNjaO4hpWOcVhJYWqxoGIPe7g
ZOnt4vfiZ8ARCNeDT4Bb51tZrDzFMKZw/nhSUJCOCDx+NPJPx1Yuj1hzYWfLLM4q
8hghgIQi52sHpn8vyB72c98UxEapUMD4HfExqEWe/dzUJF1313QJs9UxzZfq0jAx
sNZyknf2aQSrPMj1zif2ltsFCfnGIUF0gVYGkWjhJKg0Gbo545q9ubRzw/2bW9oP
8FZYhjTGQpxK45p/8B9mj1ada0wSciamd1tPAHTBYZ+ZYJ8YRownDSZJu05YqDdM
9j+BxQjSoF3+PZxFrZIszI7ZMgfrDciPRUL4Xo5yWi9kTsRFIiM26m6t6tKxh083
ENAeFLGeNClkgswmoSTwiEWdXI4uQLn+/Ay9yc452/LmNS8nMtgCYJEk/RMcZLAY
8ghUgRcGz4M4TgdswA8Fl5zcN9pzE9fuAZeZyOHNKW+HDQzqPfagX/3TC7skchMq
LImN1oTrIE0lK6Qq5qJLx2xbGiOkQhLz9IcQRZ6WxH37u7+a1ieF9Wmpld+7FLYj
/XHjQ74r7vCV5aDOiVXUWjpN01Q4dbZ+mmlc7acw3pRLw9kCKGYQx6/atDOa80kd
YS1n1llcHrZGfNtFux0+ohZNL58ZV2O+P9rhBNmIuhPiBGPVBvQcMs9pAaXchmF0
UbZlHOSObsYrium8PzCCuaop6dLMR1kBd03LCkm4hcmHxCQu5BOdJI51U1dPWMYd
zluWuALyxBe9490iAHP4nPD7YLwAjCA9lv4n0+niAu3pnxBLhXiKNcgswbyDwizl
jAe0qEsLekwi8o2J9LfopErd7qqFx57aQZjKNYMcri+gAMXCp5Yxalas1lbpQYfh
/4xprtJMdVC+4zGkteA4lnYW03GYk0Y9Y8LYneysANnRdAtoqj6qSj3gz1T2k5/J
ha/2ouE/WhnaC1Hq0WOyMnd7/1S3D/+Ys8r94/ELCJoIAp1E8vXZYl59IR6NRh2Y
TiT4vrmnv4mqCtnLz+1W/4ua2tsFPjdUtRbbPc2hcj9OwOa78EFwNLlSY97/IGSG
UbEv9Q8myESq3PtgwRJU4tCg2GpsrouRKTlsf3ES/tHCnvGfkpC0kJbGM8nKmwQR
ngaTTc0v3NASMqZYIMPEtcJJ/HHO0zlswgCKxqSwCTnAzCOmyiQ2blq8qYjP0aWA
jOhtMoGamu/Dc7KnNRj4igVBU6VKqyzmsxMbA/0/UpxTlhg+RpNlfgAtZaqckqUw
YsCHfvCP+ONWAeBKp4x5KSIr6dwuOSXldhe6BESU7x1zwDqAhv44g/gx+pmoIeKI
mIJEXQcC+HmoCHnHyrfkkf0rGNnfL6emvP4PXUR683wJ7e0Urri+ah+zUnhA+NYF
CqPsgwIRNcBHq949H+N0nrcCsGHumu7vXtPcvoTqmY4BdqnY/336wCAFoSUhubYm
q9w+MEeHsZNIDOwqcvfpdrlk4OLxjy/wKh+PaXl9PH0068bYPNa/LhWJ3o6GNVQ7
edsXbFNviHvJquceZAKKGUY3Xju4LQLXYcm6L9YqQDvhHm5GvXx8jeelpGblm6YD
8Wa38YeoR5Gw4jRd02dx1YDXPLATerqu19fGAoopaBCiMI87JcV/lu1ZeadziLxC
RS1ds4SgjuKWnS5DYDsfkek5bGaTKH3KElSUIzcGTC7XrzmT+liFpRNAUc9Ui2yP
6tcK/bLLseQQX3NETefDG+/cwQYdWNf0br0GVtcst3EQN8qdN1joAPIih+5YGfSj
t8t2OCdBjVFYhJZzXaXYs8wNOWXgcsfZuVFat0kDLeR93v6R0V2fyjQMAZtstEFE
KfxCSkK02wYbfXi9nBrIdqL0LMBWswVrGLIEOWcOF+i0i5Jf07LHZ0R+NF1WDeAr
qiT0SbWwaPtmQ4E7zNXjYToZJ3eTd9t2oLoMonQGra/YpxOeD9PdJqjF3IStLX0G
d2ZGrdVHTwqWSVh5iOnBllZEawFJWRCH7O3cfdnxb4JWwAmUXtjNKUSVA/G9NPKt
SMS8/yq3N9DufEvlM7uL+B/GtfVqHt3WhB6gnNCMz1I49l+Cm2MEc6e1kdnqc1V9
iTiLMWOwEdfcyiNzH/rMhMXZc3FGegK+f67EzZL6Df2+eMPBctDpmqvPzo0NULo8
Hw09CWWngNh58xwuDpczjy0qkgD2yd9FHwJuHslLrFUKj8AbGKOx0y3zVLgRO3Zp
xUsy0J7DK9Smik3mZ78XBZIwdeUWwE1c6hqt3uo2xKjccCNAv4nw8g+Gv6AqNbgU
y//gCcQcDPjVjBSmZdTWxAtxvyALYmeo3VozYi2xtM/mU8IC5jsXx8LNfTXUVu24
BgMR7ifFdgmcLPGKJXib2DeTioziaHOb+P7lPcePfjgjn03QhAecu97B+OXYwRhc
eiSg5VQIwxpThhr0J1uW+9rVLjXzNAo6qnYjRlBClaxz8KPZN3ni+v5VKqcVp20K
DEpkZxL/Evva9PV9MOe/ak+Fcmk2Gbyv8KPzu1sPwy+blwf81ukbmR6RSGiX8SUM
eIVJj/BBieLOFmePmFR5XM2SRWoGdjuPhNHeisf+e8AK7wH2StzgzMwRhiz3xEPH
ogo+Uq4ynlU8QgOp7aJq0vKD8UMAwZh5G/4MLwBXV0iWQzzmlw1cqWf0soUW0Y9Z
N02grjeROiiV89Y0FV9hSiNspMbIC11cOs+4HP0NRWKE7+AcdaE6GmDy47gfhOab
6mlOplbw/pv92JuV8zBn8FpelS/bzjdZLS4vO96afM+e4Ce+tUhRL1L6uOa8YRgD
sodZzZut9qjPyreP/tYvWNwGSLwi/IchFkqcjlbmoTQMo4LrniIPkOamLitKq78C
VRNotyjiRwb6q0ncPsg65SZ2eV3c8AVHoDupx4MOzv1Uif4D0BlZ96FPEeWrcxk/
szVavUD7BdcJoOR/cT4JHawOmHKdi6IeaWRzXUDdBG3AntaEt81oG/Mkk9McFfuB
mw94l6fZzGa3HZ9FktVzSAlK34lrhILsDA3am/FazXiJm0HSCNp0z14xfqrqKBx8
AS20lU83xmviILNWw+42wVmj9HUHGrOmRxEbmT3OuL1EvEOhKcJJM9XqFPyBoyA9
4OjN4zK8jkBN6yXyY3EgjHXovbp5txcmZ4y0foATUgCAWp4139/r+TwBNCKXRzrn
3WcERXFEOeVNgnYYKqt0JEKioKK+9iklCFYU0dY0mYwlpabK7lINnUvvzXka/8PK
puaPuaj1EwNkJpRshW28JNVPZ03q19Lpn2NeNrOMHNcUaghRf8KR5h0BNQW89hOW
MNrtu9K+AicfLC1fkmdK78COXjzVu6kaqb4wxP5H55ElH7bCUsHDPsRd2+84o4qr
ur4AsbEwwNCFR7/6YQBLIE7nE0url1XR0RINENk9/3IaGt+ZBh1tIUjeSPC2kYr8
KIetIrR+mp/rfMqucOgTlkffMgElgCyt68BWPA+MpnLdnIdN8cEO7wLwtm2fp6OT
GUriZCDr6rFLCHvKhtlDoemo8FVkxf4bXyy/bl64huKpgezq6dbFqshVzbyYtDeY
Wj+VzHqdv3kPe5vs9Lh8r470i1WvLTCv8N3QQDO+ebaqwwFflVdXMcrXXhOqfJ49
w21Wzs8ujWIxPuyzcPa9W7dZQ2ZS0TrHv943OJt8Uo6eTUvHXhjiBPLsEIl4Aune
Uq7bFOXdlAL6JnsMA0sIGRY4TcZWClj3ZePYcEZ5u5eG3+DTcMCTjmLbS/wDAHxo
hYEgkcBOojA6NUJ1pwYGeMgxEjLEBHCh3btQnYNr025tPqDw4I4Qbhs10FsxrBFv
hI0wyVh/mWN2Xrn0W07XGLQ4Qw2PWtfrPP7GaMjOfHZPDOV3F8nUfHKzQdo6Emwv
OtyYT25jmSX1U2rHBi+2XOMgOlegE/0a9bmVyfgSkl3kvBSMr1zfUZ6fEuhPjgR7
F+9TGdBB/hYRL8j653yYcyDeEyl4feUEhtplEisJUB6tsn2EuL7QJNKFA/5t0uhY
FgL1eDBCv83lUCy8pq5MtZcCdNHOq3ITbUeH6k9TrhTSEVVXnIHMc7+r6JR/DoB3
3c009KMy3Z+jLlSXUyV94WMn/8rVWws7ihPkoR5rqkmZUh5MYhX/RF6S/4+4lam1
paYRzj2Gz7FMI0pso1n8D5OGTJJNodRw1AV79GFlDIWtH/F3jrcSK3Q6e55H4Ycw
qo4j0MZJGckquKjWAVaZr5wy4P0FECtUekbY7fbESgDtJT3DnERhFs1IOXVyzAEP
xU+Y566nnGOA3JYflHqkW7NsF4/ES+t/uFvuos6YEJtc8jW0JDi7EMIrfyIszI2h
L9hcA0+adnxjag3d7ZYC3B+vqAfEK/gMPmdwAnrkr5tA0NWaiKFch3phGc0wIZfB
VHnBZokV/6H//huo7GmgMiMv2KvclKcs1iNLDGDNYkOamrv08MjrhPQJmDfvgdsj
ogQpnqtv+UL35PTDYTm+huQZIBF5i/knN/UQKK9tGvXJFULUKtv8KbRgD6klRCfF
ofZyf1/Hhon3RKzslxoipJALUl4Vh+WSlqu5ckx8cmX0Ujf+3RoBBZ2UTY/ihdLp
/PC/pmNmHCLNMKYPcxLB/mu5z8UuzIac574ueJsyK1fJoxKQOzSLRVeLIgxpw31Y
aK9jk85B2gymP8iSR6ZyetV2ykFp/85O34/eci+NKWvqfjs3UCock6VoyDyl6B+p
t76BCo4E6dAK/wg+GhUPQwRioqNQsfC6irrX0RAxVIPehNfIxN37JQJnqF3spbRl
H8Ro5k43axh0ULfZmytURzvl+RxdcSP1B4wQ4rjcJku6HYPJxOVR3F9vv6IOtQfa
rp56zNPO8pU+lbUS6STUHWRpq513yt9kjq5OXo72eOYAf/eXxU5HdmIrxCFDLDY1
rG9GX0A6DL323LGWPLj2qR5yGOdNta2isFPyKpXEnrAUnk120RPRHahypdT0Pvog
0MCO/kPvud7BI12oWJwmK4yyO5FbhlBknsALUjB83tqfnXldb/abG0v4uYmkWwUg
C7aIa7k1llu+leTI/vrwlJPbqjEbQVOr3LAgAa0Fr90JDGz52iPEAtcaruw+xY7C
6pX9WCe6gMFETuIYJudC9sRJ2aW9I/p1k0TTA9LPS84vDlCDBOsc/jfTXUg/xGep
+yX82kf4JCilmMhvCi3TMggtJpVaKbM5wDaH6YRkW88Y03wN2pI1Fs5SvLCohR9a
Iz/mUPZXdXxGFAJBlY8wPpcxTAY/pdR08wGOW4M7ljcsu3zUi1mNooRv72tBR3Kt
qLW3dPA6QgeTH/pAO+UCFMMXDKMxE3pxp5bnVH6WTXM82AI88D1P1/gW0ZQluu5I
PnNvL/+Yy5mNB4MS4orZLN2ze2VZYarJIFW8DPMwxxKo2lKxjYLQKMNzeJI+rWpQ
c3ux3C1k02kCaxLJDFxgMub4dDnflL9NFCCw9chJA54PPa17UwCFZWOW4wz2lGtP
xyub1tOglMNv4Ifw9zoUYkHUcrSip7omRpApIrvJuw0JkgMkKqupy7xhTntQJQdC
7zV3PT6vkNqXn72Su70zf3PvnCNK3BZhRJIakiIpojg+EWZUsqSD1wK0jUI/24qb
CJtdz6HIFOy3QLb9vcR7bVf+oRYQi0oEFiwznAsXhKCOIDNrx5i1WiGyxfyB/VoB
GTJHZrp892ERDBt3mfo0HTAtFZDdL2kGtq9sa9Ohqh/5V6kcDTyKwNNJAK4z2M0/
QMCdcKqM17cyhEjp5N1JDaH0ufD1IGsSlBrAnoKP4ubr12SlmUSxSrkxZrjxiIzC
FIgwGuo2MWQ2WccihvY4r8bqowNFOLsLyZgAP7PDbPpOsNKaiNI5ONlyZ0VeUhF2
k95Dary4TQVZ/P4wK0kZI/lSD6GOlKm+xlotWhrJub22IOckod6t1TDND5xg9NeF
nuUpIeeASGn/t0wbstvd+Y4P5KKMIIsi6fOcMjKBkgwaQf7zS4Z3bm2m1+k350rE
IJEg3SDi03BPJfxvkKwB4iTUe9uHO18rxnHLVsjugeea9HprsBoXanRgMmmTGHZr
mLJGaPNZCBm/H/A02HjFAMkuNT9HFl509EgGQO9dfvyF/cbVxhZuwVwBk7LSWNZB
/+/9NN2piOTkBf90SV/o/Pk+tLprEbRHUL6ej8+P8W0sWd1gOEyPkzFP6hdt0+hu
q8dp+MejuNzJxmco5GZs2QP3trPzIgAY6mPX6Lf8Fbj87EAYk1DxKpVpYoxhbLLR
8SpvQLBgjcndv9wTB5BH4RltQoigC5S6nDfiADjKttm8PIYSyOM8bQCke0+4LqZp
LBH57McLSi0OVPL1fbHIyCzMkKZ5K4pEACMxIqGO/z9yV1fazP0IaHSZN3bZ64MR
1fzt+QXZUlbX0UMME/1kViYXFah/VurC0EUjPbl1ybXYx3c9AswjGZHrzvrij+p6
Hg4KoEIkC8+NnHC61uAjPSeSJ0W6+yQY2HYILBTWpSpqmXDwZ3dFIePqyJirttAa
082E5dCgU9NYzH2rv3oUJiyIPQkk+KjAsk/qallPXOc1GHLq0Mh1aYjvSxPdTviH
Q03lqKYTwwuAsPzrdcK51qPcZrJDkUL8yBturX5rRf5yIFp+rYXL+RngF4sCQfjd
+cOulp+zic264GOyWILEW8/Smve0GnxkXNB6xnmMHTOjLsBc9FJUrhbj/k90Rbid
j2ESZRuWnoT9HFrnCM332QY6aCY29uZjzvXkCx+93WCgdBJEchelcl8QOo5dwiE6
eMdbZvI5t7p0C2IzlBeWzAupaVegjlZNg5tpp0bmCGglvcuRlGUOvpODVX2P9g4y
4VvEoBgLg6VLeozhBPOf8Ho4Hk95h5bfRsWSQqRuVuBIBG7JkCUN24jxzHnH9ZcT
t9TYeNw1lFQCFiQ1LI6Ks0R+ErQQOy5fX37jrgfWphXcvThQRvSLrdaafmk1pyPB
QTM2EPngTmIhHsrRGfM0CBQEjq0nPXaRQN/02cZ9GrU5tvUbFHCRz3nnPHCijEVk
IaFDGPUdtJDzvgCggidGTYUqqPp/mMuK+SayDoRqMZYYYXwQj4+3BESrJA1DszMV
TUzjiyMIeTHhzoGfGuUQiFWR95xWFLj4XKh7nPdx/WSzTD5aHLJiAR3LwZlR6ngF
g1TPgxhkVjhosSvrVWqqoFgCsOCFKPxh/tO2kGmiqtt/h3YvCmmpZlJpqGdQk5Hu
6pagLSpxTgRx3Pwgmd6Xams2PDtytu2e60l5AYWdqnfInUZ23jfnuOui5v6SOe+b
JF1e39PliMDaagYA/WJ9SkOdtXOtSgALAAMREg4RnMFsRJG0uXP++HLMe07lNHtr
f1W06DY4z9u8Zz7r4IP1ZCzuYjSOxnj8YD0Og9YxFhudCbG/GQ5wY8yhgBuC8jYm
6jOSMvDtXbQhgekgwJ1nJscHDxfOTaNJjPiwBMQQpCDRpEBdXz5gmNN+RrX/2krg
GbMNG81iVckSb8w6tNV35Yx+xICioWzuwkGwOx6TSPPxazOkAQPZ6cUrRvGyUwyd
ashltcKAHrF+PqG75kMG5qQAOuDnokjIQoAGoSgh8KUicVwZlfSWquJkVIK2l5sj
T9YCPvdKQv+lnsgSdKuDvU68c25SjCNnxGy7QhDd8yivenngHukYHPbZlWXp/Xgy
atLlsHG2hWnkUliPXzavzdDrK5PmFJvausd/KTYQLZ3/ui+AjbF9DvZ3JsJi+S5u
yzfpnYhFb6/7KoOkTngwUDmu7sO12RBF5eWMKugiKrxzw3wZSjbdNsSYYM+cn1ZG
eMfP4AeKJke0/BA4E/AlzkKKzjlZBLhEAYaQJosMf7K8ghAkNGd9DfrYXwRAn27y
shyb99WnPwTkpP/Q41CfGLpR+UZwO0F+yJOfk1LynnW9e3LoMC+xHg/5lijyAlOe
MxrL584J1Fm0j47jnW1IaGYDht3OyHDyA/zLgWJjESG/6I4JMdtvWvw8Fg9RObYd
UjT9/R5+T+gXHy1S/YXnTp1m/S5JtPPkFRcdi3ioPimtENUqm1olDrynguNiWWla
wzC0erTMSBdKTx3iEzdqWsnnX+CJPQyvFEioJsk2dEC7kKJ0KeEtlnCYwqgDWi7Q
VXrVMgetGYSKKJydcNo6W+NPGF89jgLZdqK2TMEpULujxi0Du3HXdO8kggaCvF83
XPeuBWBK9mUMEB15S8DywCCm0+JIHp2Wh8naHbvFMafMnBV9dosFYb/Leohx4+Ah
PnReRUr0ufYxuUm7SFdGsTiayMBBoQYhVg0mYfcICXrhrFQ4npyrgTjFngCmAPJj
fEOOlEcjvcGX8xuCOGvKChgAskLNCwLwOiSyYwn862p2FYJUWDmgmtiJ3MwJkJlj
t9Fo2R16ahEAPdxnpZkBSzbrk1J2beLOHRBW6z1ajSzNaWwUKuOYDgCPs9REhYlj
vwpUysovFYJAdN7OqjOTHdGsHK+7vznX8PSagHetrE+Y4CAnTCs53WbHZVBWpZxL
x50nICthUStrAF7m6qkWWRoYgtZropOsi8nRXLNy2U8Srv6Sd4AmcbxdbwirepnF
Pi26mDLDovYRDDbIFNvWBY16QprD4OALmrqPlOnX17PFs/NXGGxfF2ZZ5y3gf7y4
naaHwH7aM7TghdujEJUR3PzaWYW1stJ8yxUXqLPIighGKEynPepbqY+7+jLFh/pd
dTVxC6s22+NzBVyTUezo8G7mbg3eynTRWU2bYAGy3ToYypMR0eyXsnDbVe6vokoF
d6a5Jx5MxNLar41kJWGGjKYisA12ibdqO/HtYwc0H6hlrEMNuYwJJxpWoSDv/wcm
raZNCk/U1jN8XspSBZ8z95pBsqJIk4hYm2tIV+iBwnKR0BR2S5BPova1nTg+Wqms
2FS7eKo5u1TPYtov5BGbwuVQ6/+1cGXRcrOYzdTqVZ3HiRMHF8kGwceM9fw6dBli
cRW9RzVTBsmw2cE+qiW8Fk87IQ34ce69Z8MjDepux6KZ8OxI/L9ON0GX7V0kCbFE
fokJ4qTHA/08HgY6nPXyibcqINEjoTnpT8fRrNtLA2bcEHaX/PvoTd4LHeNtuV6Y
Lxv95En9kIdltU4p8tQQC+DqQJV1SjKUIKhqLMLZAPCIAOPLDGKD7iXFVWhb0kmK
JM1/o3bZeTU9zCQBoayG0JmtOHnOGFwagzUmFgGF9tsBFtE2y5V7aUWG4uE7Jtd+
jDu2NifAVbA38wPjcBvylrVeGwgMnntxcZMQ75UJb8PN+svdIG6hoc6iQ7cuON57
znx5gRw4T4J5Pr2aAHNahfMweSE8OdxYncg2+mmKJ4mequQ06XbfrZ7JoJ7UYVRb
h+JOSl3ZzJlEnlnJrtn19fq1Ibg91HIbF6WdIXRp6r5M6RJtxzT60V8cObwPj6l9
NspmM8LLFCltkq7LDlgEaDQ1XxW2VDsqvz2qw/1+k03gCHpD/1Q44AhumJYiHXz4
R2TCHbzVVr5dwB+Wl1nCsIc62LBPlTMaEOtOO/TZ2Hk4fCL92I5ZuqPTRLZKMZN/
YyO2N9fjQN2T/8zvmgoFMQ==
`pragma protect end_protected
