// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:59 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
irnI7hE3Cop1+V89zdf9sa+UD0L7ognPOXQ2nILVCydP8tXo284isjj20qzxaPwf
YjjFe3Tfe2mm9qAdXhqgrM+2wYepera06szQEOPTe9j9CBvTGMBU46kU4HZK0Hwi
uBPM0hxFfsoBs1I2E/M7VQe9OcZ5Th2YIbuwrhWSizI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
qb/1T7K6WaarZe4rYIjhzsxPtBgAEjMwsGBCWdjCgVd5n91XgpZKUMU9QLtQy7H9
jt5tm7ezOXRGI3oB8YV9pGutEoDNRcqsPhAYQC0SjgnIipH+wTD+vs4fQqvr6Gxp
K+Q/2SF7vmDk9zKwn76FDub7SEdwYFAVVy9N59l5gxrS/kJ/uJ1UtYPNOwPUTDwN
GJu+zFRXJgKg8Ppp5m0a1L+u3a4/xjv5xJVnsJ+k3GW2cqIPhICwtKfLgtgFPDF+
Irq8drwcjwFrsEv1FgkS8jn+rMBU3u9dErfIxKDwsZMk8Xoa0p6lnSbpREHy2k8b
XkPK5Q5EW7cN4GRkqo/VFCNXC2RXktiDpOh0dLyISUMW3YLh/yC/vNTW95iK/YkJ
nfLxt1pTly1TckQz4awmhANsug04k0JNaNL2RnC+ohVhnPdnQfLsihGMXAGbuHgw
sNBa6QijyyYZy6DNlIOV3oWIKUVW2Mm3Nu1rFp2wBWdGTYKsU8mRBmbgQd3V46hx
jTEYY4ddKZ9XY9LHHNHpsjBedr+IGsMXmPJMQMXUHPxCxSnrit8p12cC8kWJrZM3
qBMX6BbTEUnllzg+/qibOn9OBSyp5DdGvU7bzcUIEaryU2kctYIv+fRQvGnoaS21
Pmv3t6z1XWZsSeu5xvjngLAkP9u9OTa8//LrX28/4pCXG1S7B98mbs1tpyjDCEdI
I5YP8ozocT/Q0AplDtkmk7/85ehSGqviszPMu3Trhy9f4jvT8+jdYq97Becp12uM
8E/lgrf/Yh+YlB4JEE99dmDS6uol1FWHv+QEEriSm3WOS6OJ86YJaMbaIHfNVZfR
XAboNTIgD7mTrIOwhJFgbC36BBSt+7vn8idbtCe/Q39o8UEpVc3Pn93KdRPKeOSU
P1ZCVuj+Vb4e1F3vio3rTZwF0VJYwx7z4OM1Z8J3zJuKxxOrgFhKOZA4ZpruYQ1y
geJc6F5zZ8xrqg7kFvZk6rPLpBSj9vfyaJnHzgOlEgYeC6bVtwvSGKN80M3KMYDG
tY8doaSaFKmhIeBDudt0CU4dWneYG3nUYoxamw2wyczw9McDPbet9E+Re1QLZsAa
8wV4Djy6V+yFvKBaYI27/AMq3XMc36dScIUkhnJ0qL9Np9HrpMZ/pRG/oEFSqJax
9/KoIU2RaQwMEICtTcaqdgq8aits+imITEki04vRpDK3qfzyTOLcsq7g0znjF35e
yMa8cr+RtaKBiZ/gMDIrHS0aCCeQl+NnKWVpudHVf6GEOwMpTTNKuRirrLYeGNLz
4Am2INabiOHBl7F43JsSPK/NDPZkY7E6yyvONv41ujZh7qXLRkSy8zZIItDfQFt4
M2eZw16bhZLi/DOl8ZuBJTBgHiHJwazymc8VvcWRffBYdfFWHv1xNVD08HqEnFDD
AAHmKnQtjO+T2Bk9liRYYa7hzURTIWX5jwhoxEWEaab0NUAmQG2UEpjFprENaBQb
R7+S2uEWhW4sx9SeqewjCebXAcjcTuuan/JWz+pDFDlHoMBu9Qlfo49rK0rYTvNM
SXc1/wcP+U5sSL1uzTnsR4bSiQ83Hw1y3gw+yVI3BGJcIj9Lgr9ONPr5f5Svlydw
Z9Wal1WlLqgNsKNlc2Q/ntBbHEFdrK6XAn7iGhJPCtfcnJR8s/B1Tu5xdWhlJCm5
Z5eGqcW1iqJnoOtqTO7bh8PyjaGpHp7sOKGQYQYJwTxID7zRX1ud2xXksdkmGG5i
E+cysPWFLFdRBOuYJUAV3+DWKMkHnXFLqqNyeA9dH+/vL4mTlxXZT286p1nh7htJ
MYjv0I/Aqst2J6sq20vaoOTG5WJJjrVVZmGK3lmlsvR97jppw+QIGKFzvZI56Heh
WhkVQkH6HqxAhiZlGIjWPA4f9y7Kb48R4yCw6tJ868AUv1QMApXJQPx1IezPQPB+
vS7X7Q+3aZJHShRlFlb8iMTEmigWJS0d6nQ5XHiRsvuIlsyHeA6OUJxEOdecwP4P
VbDOJSloEkUS5n1jhZm2ymMuZhZ/alTcMyrD5PDvrIRJfxaAI78n4JlPKdT/Iowy
VbQsmKg3KWkj/2OnPs2NbNbkqSL9enOppcgQimRk4Paddz05KXFAuyAOevQ5LLeq
IVbFUGEo6VgrW9beIvYUS+HZNKDnIWZBFmEkYjk3PBn23hbCFh2a68yj+bRJI2ek
1+hbcDTr8KSehOwl4VnaIbe89737cy2tQ0YDV1hKWwcMk94kDr0Oqex4nEDhxdMW
RFVEBzzO+R0e5AN+lZ4nr/CkuMIYdmuPd0VYb5uWnRW7vrgh9281GMTBdNHBCnNb
PDNHjg3MgWl6Vst4iCGNfPdsrzFa8ikXxIDU2UnFdenODnFVhhVTz5qXepVvfEm/
73x4r3U6E99fkTuCd0o3Jg0KcyauL7JuRyxji4aNICSl7JP1mm2p6sC8Lv/VFs+t
nJeoxD/KkngsoENxjMNtHTxVPqPAUg4t1EViBl2TOsHaIwBVNwnuv4Uz0j5ccuxW
lUbLrG6mk+EVbx7IB2zzOwo6hFD1iRVDLsSqMNk6LWmrHRsO9aGsOJSTBqBqocOn
uo61hEIcWLbOCoS3iRkxr90lxHnu1udrMKKa4w3KiZTzB6MnFfoNkGKp47SfErNJ
JfOJsMfKMMn5FNktYoB+SlZD0x2Cc11CjB/NE6bJCsWUU8Aiw+H/bofntlpjONc4
rWO985EJ/qdbwY1u4E2Bmz+dVAiLIgoBEpXiMM0Gz1QXMLBOZ9wqrqENV0rt9Uac
4Ymvs3lwAg4lHSAXwFwloT/WuO+/Rdk0B9WP2KxoCIGg1Rks1B9DFwVCPW9eFmmV
xyYZpZhnfm/5u36EHamOU1D+iYvVjQLsjGjeokd1o0DVcQ/QrLZjZV/wTpSXMA71
C2ViyJWnLnTb7NQlrIGad0yc7OOwajoKWnEXRswk/d9ga01Ftm4JoME7/pHi/Cld
bxnvWQiHlqMbpWrgfEXWUg==
`pragma protect end_protected
