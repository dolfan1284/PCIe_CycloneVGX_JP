// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:58 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TKpEFKHBeOV2IRoY3tiYbeukwHeKEJKZm7v1tYc7dDTYrxYTy4JRdGrlkKS56r8z
1QpdxRYacIfmRBUEy6ujXIgbTBZ7keEgeN+kVs5JrXaOs823hU3KsKbxpx23Onz9
Ytpjjk2/vG60evs4Z9q74Z+FqtVcLnlOvmDgQ6Qlsis=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
eGqoD5ri+vBkenuPS3EP7k7igOpZWmia6JI6ipofn0OK5IQo+0cUjzlgsFhWTHBz
sH0ncEjOqf99rBi8z9mstv4Rt1amAN3de6G3FCXx4n6HRE2eA1uvdlWhKPZ6tqcz
JDZeIeYT+nt3FrdBRLbVZQUujmwoXJkKhgplq34yH0rPvNLGbDCxuUvc1jaNns1G
Rtxnz7Lss9uOWx/M2pgGjJ+1PN3eBcT74bEGC4OCliVYd4kZ+7F3OgBWVwx7BN5C
keZg5bJKN9W4QYtFjHk2yFQ9UoXYARnJI7LcfU4NiZz7JvtRaaGRKYLeKUb/ShFV
0TKHPimVrsJRyWt7eiYgNjJ9n3K3OS5KKnoLACyGg+3gGbK6LfsgfeqNpYPX0Rg7
Xiz3uJSwvn0+3GeMkz8OU9penu/oE9pJam2Vy9/Qv5CG66EkLWK28QcyLTsmnFMl
u0/EGcH8W4Qn7+8pUF3b+pM0uqBYRWxk4zvjnBZsk1RdsjdndKBIJFBGs2V9zi/j
xvcZ5lsXSkp9a5Jh/HziQGWsnkMZDV4c2gj6q6XgCqDSiXehZs6+mqEGq7enokFK
FUO1eM8RdzZv6JDhLnSBVYvQq0rG7ZC7+hb8eTcUxEmYXB3na8GGMaggfZ4O9I9X
BUnK52WkjavSB7Ot8lpO9MjHoBjxiXDMzHUQhgdmmX9CxlHiI686PsQlQN2W4KlV
XizW+MN40851a5VpQbmPGsvucEsMsq512HPhar8wgvtqhRvDRFMYiONHmuGKhnOI
i6u3qxBoznWme/v37I+YYoJzT0dmkhkHMJkZAmQYo0pq4pCApJ3b8haNFwmXXamT
T3bOG0DvfdRmaVIKS56CSXMXYtpzQwNvJvH9xU2ED5HDeq6JjoeFKOlNlDtaoPbq
o1OyWRTjp2u6hpHxGR3RiUGko9Ek34ARaG8M/KnnSz+no7Onu8hoC8k4uClsSclo
CpX14FMldD1UejkxsXNGqtM+8DUws+JbOnRT3ihiZwv50isV+Qhaompw+u/i0kLI
2Wc8eP3iYSEM5V1tfXVEaHTPY394QZ9LCJIRNXoWQ/cahm6UUUnp1MhYAcpJ85NP
JDhYKKxFkhdPCbFmNtqZitSkPvrtMbVhautIqlLnNsJ3wivvejGP6K914Gptffoc
BeL+zCc3fpSvnqKBgWcVwxYOllnDn+SsYJxdFmKVnTunvgWImBJLy+oEDFL5oLoS
S845IjtPvGFqQCOkELVNlaGpQW3+oTyVtUPkBeL/fKu6AgnwEMt+QFdPf4u1t7Pm
PUQloudOQI98Tces70W1Eyeu/sG9PHFwB9gPAQqjClfdeuQ0w4W8xo3IJ4KBRZTS
FqpxAasa+QYFMdoT7rQ7FqAZVpYD7a+Bc7yfygqQzc7Fpd/k9PNQb6Mc8KoNRnx0
Lmcg8vnp+h0v3npYQL2say50op9iiupJBNTYKwDMvEYM8msr5j0ph7SGF93vfMa+
myndpQn7QcrD9rjW0IDJrJDG/PupsKpT1S1kcGVmZgCjTDscmcaNRpkekcXjyyrl
s1d+xfnYoIbBrKgkT2pCrDG65raG+QPYTda/h4g9Oh1B01XfPASzGvSj2Grdi2M/
6UFtte2Xn4UvezrZJfWijGjyPdVf1TKhG/3qYhpK8iq6prENnk1WFAxOJOgNeg+f
OeteAW/5xh3zT5kgr+8kSVnrHTUue6coOBnnlZRypkbPqGm0JW30UxrHTveLvchO
cJSh46Zzsk6hDiw1AcbNHW0Bgr84IXTJwAidDjW1B7BdhjWHs3viImjAcdSH5YWj
LMJ/L4dFEGXJ/ujoU9P57IdvHOJnthC2GtsF0BlBRMlduGzeNsdY0dTURHVCAtP1
oxbHs1nutohlj/sDow8irbLbTpR2WUO0XHvvBjaCl+ZhlGnjcyiF/nyxMGQpAM+r
L0q2Oxv7FYlkg9ddVnglwcS0dYAZLDkhrZtFVB8kTaJV0jReIY6nDcUWzuT2rtXl
iILXuUOUdWjZhpngoL2iYpptyCXzL96R1KHSdaqZx+RfetbfZay+SzDN8qPOTYZI
2w+x/b9OWW6eC4ZVVAImCRXTj+MgDdxitUx9pOz+ONYpW5QgYy4xu0Pd1YD6WB+a
O27hQFuRuS/yqMNsubnL8Z0U3lL6gwpb4f0/PD8bHzWnACofTqck+KCNt8MPo6W5
EXP3LBNzTqVM9qnmdQJ/1lxqQT+F7GzqHnFNC3z/nJYd8cbavpgjXnJZ7HVU31tr
t3L/1VnItquXNMB/2klNswXUuUx3XyYJAqzyO/fgaV6aN6dbyo4S4SDdoNRVRmRA
Muz+0cyhnLb3LZo9/gx2B+KYYJcH3Tca9d8jp7/MCkLZsZQuBeX5lp9CnYQyWggy
KMbON3FO86TsE9bZ3r89S3F5t/TJsdiMeD4aKp/DH8Q3TMdlkSf1BR8Si5TOo6UW
Ky+Ae1le2u1FbD/ih43r2AgPbsah22LeKN9BkmOYYkcnARMkVYEi2c4jAsorWrF4
ypH9dXFBSwDgUUV9hJSGqpyAuHWQQbYm6/ewq3Y+1FgS0pkJZwAB84pMdovW+oMm
KDy3ioDBpfY5lp4OQBWvtMDds56qm4sCBbr7jlXzVOK5U05Gzxzv2BIICfG1PrGV
SyyyizhrvYJSShjX19AnonmgmlKT7iKHeOY7k+9W6vYJKjvDYcKIXlIE54m0frE5
XkN7OJcUua3+o8Vh2P2gJ0ruwz8HFAM7hlhnuubziNoH1ot9jK28KqqFNvStuzv7
+b6lasv8vvoNaUIUDqe0/vhRO86WsahL5rlJRrnj7D4OLyJGxsJj7FnYcpcoDeuh
TgFbpDYUJcCR6INPTU+k2wAlqxOMveINzJQJJXn9btPz9dZTOVrP+q0XWCHC1KQf
VpOpMh/zEWw93gwT50klx00VKwTDQVGA451zfvFu1R8oCAwhzo17RLusX+jD8N/t
KLSQxdw+AxosuYZ1IAnvENL1DKIN+kQgtI7pCVW4hgd8Ub/uzHd0OqsdHytfe4lf
9uBUCu67ZWyFjnIEUmhsRJg1n9Em6p+CKIpVLKqBt1fJcsmxTqwKuPd1mv4B8xfN
i+et34cCTqgpHl51FsCRfcOoX2VRsfCPX3lpYBkd8DowivQFpvgZMP5S+ORyZkCB
9QCOJyDO7Vj9JR/A0MpZEzbewj1UZ4lPe5eD4/qdKyzOAiwFvpI35Og23X5dnQog
aUN5r+t2ZrXGJTwQvY3Uqh0hvwk6lgs+C+E+r5+9hXN1k8iDt6Tn5qIBBxRM8kpq
HGcQu3rbdgLy1A5LjopVwKfOZij+6aw1AZ2RqHF1Rl6nL/IQEjScxWTOQ+9EbtD2
3hzpF1L+7Ez6SO6vABvWTnXhgUtWfaRxNApcJxkitpsVzQn4XTJmNuc1q4Zp4hrw
7JF+PbFFNvXN5+FAd4u1fgtWQuafdBtQxkkDx0ruXd96LaDh4RcuuE0NLRKxuEH+
IAK8cDd2hEVo78opDW0Rgcj0/fTEkuAzXQj53uDdnWAGM2L2iWqrko5mBBv41GgE
6iF2sXsG8neTlc4bIR0wnLNeU+223W10HwUpWOvPWDCuWMxMcm6wQqdg5QyDc0d2
ToYASpWs3WrWY50pg6eFAER4GAGu102AoQ7zCSfvt8+gxYYRFB9CyI0grPN4Ueuv
mCElU8TcCb3aH+q0ZgNG95x8PtGlXWvoC9RFwS7RLwbbHLhu/lJ2jA2qF5aOAWLl
1QZg6NLPyqydqZo93q1lGm2ky2jBHJkzfMB8n4P3NubXM+gCNFAcZNosygZlCouo
wUqaSu8m7UR1pxJK6U1QuuU3+bpu6s3XG8bC7g6xNez+mWQP45F/wQMxDkLRT825
aVV8wrLNM3qnSdj7HUDj0AHl9SPQf2OV//20tf1S1lJRMUHnGL1NxsbUmvOAWbdD
yXVz540ItanWDp/RmZZWntrPeetZe96FTUZE0vsjSXxJ5OF4p4v4X5ONWfqNoor6
E5o5zMY5f31lwnysnZ9mPmUaM02OR7T8C1KfHUJG95ItUhqTUZfqmeFFMVWP+sGf
r1HlH2WCkBB1vgLWSEiGi2adCDJYGkczT4iy7MxccajGRx67s6aTC8M7vcjxQjDd
f9qA5p62NcXaunb9WHcwMi/tG4ezF9Kybb4GNYFgnFrbfsEEyamDG/2vzOwdxTE+
AuzE0syi58z+VkSNZdQA2vgxOnPN9w/oeENB+Y8sG+5KyXQuxxAstSDtx05PpGYu
Q6ylYv34oMPqz4nZmCTUmX714aQ86iABsuQz/QW9LqfhGcG2tOxTo0x4zLb+RESo
kZ6Zl3dldBmOLNE8eAbguYIJRgzB2DJmpw1x7cd96xYZEQX8O/JtX5tyos/z9kfK
/3TG8pNboLTpEuEiZtbI7ZVBgAsCKcRkDV2hAfGpZ6EIyCAjvsBKe4r3xfaGjQFi
fYycH/GDEeHYebPxAlZStWENgsyv8Mh2ys6HeqNR7ywXNX/6w0PdrA5aSGbUayX0
1raTBOnu939Yu2AxDtspRyZE7rq5diJNWziFnWklJEJ7m+ZIOONuJ1eG22RWu0Qs
dBxfabEhZP85P6hHN6u1xJjf0iEDO1ox8FUUx85BrPQkBZssKC53oACb6VGR2XBA
Qb3/nFbP0ypD7+aR8GMvag/8CSQu8HckQVYouXG9VSTfKwWWF2dJpoqKVOP4plup
xCrrCol47Oc8dZ8uphNunHA6Tq0lglm8BcMbqCf8BgC6ZPEEWraGWbD92763J6Pb
M5wEgYHLZpZvmz33qzsYNfJtef18Za0BY3JKnf5EOhkcxLUOlAiRZUMz/3uFIRkb
QiShvCgIFq6y7lWYmAbcyZyDW4RqgIyRVXYz4Wul7Nd4Cx6RGL1OKGPDBC6YwvGy
i8Gs0sfGT2cMklsCgXD8cMCjauPwuazwYM9/KzUVLeH6YCU/Rhi00Hd69bJ79lTH
yMEdRh1pipw+r9khg4gaUaLn4a6valLnLMwL9dgmnii6hYfmSH2mlAJkVEBFU07X
GHUKQY/In4DQy5LVJOR/MuG5tLRVmfHbDRDZxGNeofV0l74MGNbpF5O/qI+DDZIa
5ppqGfDzVy9lAm94Jy/621mnwnDF2KPDLzj9KhdOUXt8p0blkZfKN8tfBe8THwEQ
rJ1wcxx791LmsU7LLFTfuoRr4g/s2hVLY7eNJiQpCyTDZu6P00MjrLuuSkmpn/RO
4tmJ0jHxywtdZYB+MnNSNz+jyzgMAhkTFNZeHh9HPoNfIfhcgeUhKPZ5Gdj6bQ1T
j9JHUTJtm423NfRwZNcv96Qv/42gDYRi0Mh1q4CPJpWIXQB4wGiPfFRU6Xc6Zh8V
eQym2aVNdDRbwkrJzG5MJWhmbOzqE8YpFXv8JhasIf8DJKS9Ve6eJjzUKfEWFsWp
TVX1M7Iq4t5nil25YlKFOabvoIKvZIp9k07cznaCRtBil3nIEJnOze8SzvqzyTzu
ZfiYar1SHflozCumYlx01UO7ePLE7u04uo1gGhnKA1KGIwvIz+LUuEaHhCRSkJvz
1chspGuWUPh3Bpq9GY1GFuYXKshfFZ5mDzptKzKo9Fr3hgfFgj4mKtVnt/c03wV8
wCSAboE5DAcNeyMWVgwoHSxtWVeRJ8KG2L20tpRb7fIOQavmn6A70uACneGa61hm
GzYeKro6UyO58JzY87+XG+mrNCJocvzxBvRePujLgRivRksWnqlj+rPX0LFzLE2s
LMN2CWMt/1nOFEGVd0Q4Q2w7JlkAR9CQMmpcnZbm8JWK7Eh7YRLdF7QxeahVcOOm
cD7RHZVSFvERSY23AA/e3cAF+8JnC/Fu34XIV8eAXYF9WX7fKHqYKmLgKf0jDTqL
ALjzaaF4ZiTXTy6+LvBsHEuj0i+dO/Awjfbzu9SaSdLCtnvYdIXUGq/1/5x0mCQo
Lq7MmSjX6x5bCV0KQ0Wymo9u0wxfnQVxaV4JK9TMoOWd5eMq5dmJp6ZddsO1dFse
ukoBl6YAk9QFFrPFM4955GsZ1kpw6Duqm+FyHb/Qf59vD0tBEmPL5QkIBinH24zb
hxhf37A8Y3D3ZPaRUd+HhmsPBBDKLFoO0k1/31uDTj8VGgvRi4fLX++LDI9G4K3W
eBmuer62Ej+xKUibIlPw8K9lvZwLnYFYxFhCtJQLrXcve9VUh29ODRRDZ1VJM4aY
IsinTPZXDe6L62PdN4EF9Uu0UfolD3kQlwMn7FZMWDC7sGNlDazvxQdGxbRL/wRI
f0jg4B8oxwsDhkflYs5GJV7CatcKByhEIJUhCQO3jiuH6O73/keEzQ3hoM002apn
Vg4NzfGVtffKanDMP/+B4CtbxlyeCsmgFjGlGlxm6HRrWFP+p60/lQWTPJSKb3Vn
twrSNAY8MFNd/0YxGoYuhl8XHJfgb/OPLDP8wmjDmn0xz9isYR6qNqftooXW8ZOP
Oe3eqQuSXtBoltn/4eWQipgKmnwOpF1HJ7N6zq2GxcFNEFTye9oxk3VN2ksuHQIH
F9UvfFN2qpEX9wOKmzObHK6BEUhNoFFttHRDD3+SXQyUVVWq73sMbjQQDUQ/f42w
udEz9FUd6hyAGn0KHer7nWb93URmOk5XcEUNELtL64rIAdtwklGIh8ijIRI+BD7A
v/XixWQ4CUKNmaRvFUxr8rcj+zqFUGQpnkWdX7jHOZ6qR1QlkqzTQO4/iGgLCfy/
qZoWvChsR9iPJLulhGsDYt9KBjDkhx7of87fs24xyLq3O4E0AmAWgqfonxeyWU+E
yFelM+iA+FDnDEWCNlhArtC5zMo911eVHo6CKSLT+LvOkyih94UF13bZGnbXR8NV
DTbnvF7ZzLthe8qQgUQOLmIfwXGdqk3uIvfxTSsqC4IisUjcvge5+TJTdvTePd2V
rfOurjnIzWCZjDpdaa4GN2+WFQ6t7Z85Qehi5MEZQ1nteWgT9cgbzoNYDHKU/he4
NPrT06oMsUBjxHNjuhArVNNGEeULFUWbdvhdu8u/IPLnX5DCvqYWPbt5yxh0i3O0
Y00J37UWUwn47yCqZWaLOLaBwKGFRuxBgqCQRBB/7r7E5L55fmv6PyU1AnfL9mj5
0/olz8bbZMOp/baHJimiRkif75dn/OhI3oNKlefLA5D2zuMUJGopF8nxr7UfN9Rc
NrXMcu/Xpnf8+nYO8FfD1D5c16Jfv9jCxWLxaBvGK2uLQRyC/xDHNzZCn0laV50L
MjrODIxOTUEAp/21jWaRTqlaqBBrO1nWYuMAGiJH4QDmCY6i1f0nS9S2JWZG/KxQ
QbAAN1GktOduU7QOUtyvt+R8VPqlJbSNm5e4D29JHJw+Rjoz7jnyH35582aaREfl
BOgEEteEpwIYPJgFubNKdTgT9jOeYpd30j6fwNJaTXaeAzj9bWPiDpWp6y7ULxmD
RFwpIZRKCpINPYssKPRr7wHJ8FjfVGUtH3mladDCuogSrF3d2vsQ1eWw5xn3imLV
FKb+ZbN8164MPIXVsd1ETAcZUsipQlHU9vVbYuI5Bfzxel3F5NYaLherp7gfLDo+
3R26wTtIyyA79l0EJj59ZjXIlPY78azeQ1yi/mcNcgtsSrxoQS2CUP3B/Tj54fe4
OpO5Qn8mR4Ovn0YF4UahfYMnHVTcrbFPCaZizF8w46Mb78aEA3nifKNzp9weu/OT
vABZAg6mYfgyMyP+/WceTo+VC7Oa++nzc5VvPOw4+P5Otjh6nGXjayTIyTinYQe7
Nqit33HNo3Yrlkm1l9eqeiZP776dXANPiZsXJ6yOge12ywWdbCYDLHV+ygr72ZS9
2fM0/2ng5df5IcZ4o3sgVrdS+3Ss58EXHkmWhPET9Ns3AUzwWuJEf4y+9Pl3CrZH
6WAWrxPmVHxZxU3reT7UA8aw8E2m9oenMVPJ+f82MRgxV95SgvitZCVEqcuV+I/X
rezLPgfBYvFMbOVS/TSOIRPr3gYt/kd5CLu5iXWRVwxkRB3D9zATtZICiTYe4gSD
0tcSacFSD/QBtmR7HuopDooLDMb4Qgi6npNFpRmJ5y/EK48lEzrypRvEymkGNtw7
j1lxDFPNkJcoBLcWf1vE8ywZj26eT2sWsqtBL1sSQeXpwA1bNn3orEn4P/2Gy+bx
JZh2n0N4YUc7GFR20dqHC/k6gms/Y4FwygCTYJWv5R4KfUSnc///8jiu12MYX/rc
AchsQETuDCVR2eQFOzKjXel6Vo2EcKcUrcLhRB4mZvtrOnm9GAmEndLNc3R7jxfa
EB/K/c64l3a1MWpFHuGtNzRRvfL6nQKFVQDN4v0vuPMzXRWXjXUQad5wlvw84tw1
TeDW3gi4OD8mBZetd/R3xNitXw8S8eKqztn7ahdRnHNZ1gNu++SwNM1k2LZzeRAq
iGxvUjrz+abvjCdYYpgwehg3PkuCXhP82sYf9PMH7Q4LFOArjXJKH35hWT76QK7k
dmCoBA97A3Ez0nTuuunIf5MgXjIN1HuoT+ZLKDDONp/hKK4IRJBZ2W6bkayQoi+6
BZVO5G5ySRLhM/LRXtj3JShiWQITteiiVwJqUSJyCUAWdXpxL164qJPPnZsF3AG9
WcmrzKYGgyOyAu31a5IVHanX8p1o4VRHbZiVm0Rvz6YEI6SU86NeEfeVpbqnWV79
6GJh+AiHdNF44gwehsSyAAnSTv4H+ytBA9XFShjzoiTS5z6bTjjs4hQI+q6GWXDy
Kzt80Da1lkdgW/vjm3NX0moZXEqgY4ao8oS27cZH5cbQ/W2ywjLPVlbpY0tl224p
j2X+XZnjXe8cXzGeKwRtcD/Z4jS5q/UTy1Z1Ll14Du8J3ZC3MvOZm632FozYrTUA
sR2ZqLxFcs61en3UYMvdmTulSbG9NdwVaMvM1MRQd8CyzaJXXcLP1Ez2uf8PWSIw
FC21u1YDhp0wF4wdF/DBbFkNNH94fE9OAsWjd5m3ye/dgEZwz7xThQODfiAudlkZ
BPGUdZ0UXdb0PL6EeOHz547JA/bx9PqI57E9dA7wygE/bLQyCijQj0FQQ5H2mJf9
XiSx6HZzdpLMbbbrMicpKsWnQb2ISPilPMRMKqD2GpuhBmy1BhK7t6BNZpMHvTsY
tQ7MHdO96aArcv0TXc1qkvyN0OBu3g4Dw+2RDE2P3aiz81qopaVk2ME2HLrKmpMY
jdiYZqlziemMhzdWWJ/XRrWbhNJrTE7BFdmi9DfHl4Sr7zkNUfFLKHEhgpvSWWYD
N7AXDMqdLHTJXf4Z8Gr2/y4H7Ce2RUVp7nzJdA/IQtf0+DezPni6M1F05vPkFpo9
9vMV9v+9Bh063aOud5SZ4oub3X1orIUgBR4lw/fKRTOZdgpebUoIOUA1TMJtRi+2
d7AmLQXttptGgXRqxaJs9O4M0mPsPhpKthYAwUlgVFTEJIpXqOkANh4bPUy1B6M8
ZHRDILFR2yU5TYgga8HT7hGnqtltm12oKLDEU2Jv8isMCsGpBwKLAeh8kUV1X0jq
FrQn5SEWuveUx9udGv68en/97gJ77gJWjHdU9wLGzkGFuKPk87gK5a0G/0cdQl9l
dow+hChGGkZxAfeGJ2gf8Q+T0Pjg+sPtgtMgHFNY5w8eirbvVE78URz6nbtS4udw
ZHu14exyFi2xdjc6T9OyfsqK6s/zmXq7DUz5czE4v/hKnGx3MPa8dbhQ7coxhl7B
dX1NnuS0rCICq+OerNQz2PQErZKNFyr3mEQJ6oaMVsucVOrqo5Vx+iWPqerRlU3V
5QgiDx7+to6Mhr19qX+uRiNjAwoJn5HRHAnfj5hznrb4bEVs/Fk8Hweo40jrUs6C
qu3Ni/YvFKOkz0ecS5N2Jp3yU32nhbHgehV7T+A9UFLSQs6RgnNYF3A5fWNVs8a9
kY+97Ty3Bj9Cjsr8vXXCubaNPWroSkdigYTje1cbn5bk/nl58O0nbLJ5g4fnWMza
CPBhDCFBulQcCZZQmTnO4Y/SV50J+CXr5xJISZh0GvNDaAHyJ8VKAB0jONY1urL7
CMsi/vjYaRupJ5vMLbSxg7y9xAT0PFBcZzkEx8NR5EQScwABrwI7PWsxqFFg8yqA
0Qpkrq7ZJ4fpCgMo8Zq21Rf+awd/92ah380XcufYMI6ZpneGwKsC0p6aEXeIo6+b
SxuPjxhpR22v261ENyciHLmCTcCo+LlwGToEPLDAj5vD+dZlcx7IuR1fr+lGFK9O
xScVC6xV+vJKoTkWHBuS7QaxfpH5sJwhT2hQBrWAo88qCShJGgGsr+bW1Mg3w2s1
Z7qWz4sp3lOW/Ng2scO53eP+p4Flk3xvIGPAEEauTPOh0WBO6ZwQ5hWOUVf1R8vv
qIr6wdr9WG9AR55xEczte4XI7S5ODvvCmiBkMCcxqKpSyKysfREe8Boq7L5kA0LV
/ctC120LYmlIcUFtHjIDqiJLllD3Gu8Z1HAOdVxOTQIw2/RJeAZwJRS/P2UaKFbV
Z0bYOVXrvz13YBWmBQRlOqzYUQl94w4hKNbAWTGQ+0Hn99H1caz2sNOv0OFvvtp3
OFzIAINOmoaPdfT6N9WGqFOcgVUwxYo0LDtC+A9BzdKP9q8YIdwRIDJiPreW+Hst
IBrDLkmdMAJTUZgBXyIxIVz0x840ZNMl5KtpvLIbEQ6EX9dqk8lsHctkqGm8i0db
zpl3x+BkOnOr7OMuZAqHVUW84Z+hzbmvDF743M5uaSyvC7CIYKt/JyexxTWXP35p
fMR1x+JCUeVGBm9JZ+54l8KuLtFjWKCdvGQPklwntnTiTMykHtgWuzBtIRwW/hl0
sOsjS1b8UXTbhrUeaTcHYOmz4VIaDI1uRUmVT/XI5osIuFVC5bYziaejNYoRe0Pz
gd0pZby2UQaIZcLUTY/aQKFUkXrM9lodp0flt9gWKhprTYmIrlumPcWMxcHwsSRw
GHqI0zno8LLvCCW/I8oyllh/LoD0cCDAOKbbtiQTR40=
`pragma protect end_protected
