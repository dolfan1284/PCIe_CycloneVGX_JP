// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:36:56 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y8ziEhzZ/xSH2ENUeDWulTPpZHmBHH8Q0qxG32aqX9ZN85m7SUPZfZiRH9Eaycfl
ZWLLiLODvpJjrDMsetmOmiKKrJkKnmo9kO10n3RzmcD7SAFURq37Vx0bqxieBJWf
MKZcW3xV+nJu37s4GIoSkxtltFgEFmcmniNsWzRJ7QI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
s0UvPmjfs8pxz7vRf+9e9cdBfoqebq30VkxeeoOttKeFUIZLtMpt8gerkffjoNCH
Pb+MT/ncUaUzvsSnaip4iNrfs2oBG3X8Sa2/nKaS63p2Y8HOIhrrdtqWtRvXB/dv
+D3bitcj3iC93FIAjPWEzlZN0oHbBSQ3s6WGlbSkKUUvTqEl/99o1EmN+Cfu3CXv
SunsGXM49nLAD0B/wKRIgZpttcCjf44rygA7JSV0objbNVzNUueeg92qkG4Q3cNw
NXD3ho7Kub20Za/g57JswqrUpiP+wcw4Dn7G8OSf9ryzv8Qw7vXLb95bRz3/5gMz
IQJQ5AKKuunOjxvWas7ciCHWIPZhaEvIGpshZfB37mAtknuqNmfoY+qgRTCVJFaS
mnQvXY9CR6iX46P2Hf4lPzURB7ZU5hW4gp2UJy51t/d27Y+jETvK1hXO5kWDngV4
R5yyBeueB2V+qUEfc85T4T7Ert8tWBtZcF4sQx7jaBWoatDkHk4R8CNvj1e/uxba
dJW03gTVKG8aZFXlgpsqCq66CeKV8cvLxRxrd+GDJtCYrnVAPzitqbIpUqqA3zbI
L23Zi272MiwISSUpLfGu3TlNLYiZRW4dQBEfu2W5+ga/mgatcZdjaGHaVS++b3l6
08z2ghiYDVdZWM/6U1tq3PS78bNKwdK3LMw7noCKzIkGq+kHnIxdskGRQVtF9hUK
ART5TArTwBHimGzjhcTSlV5z4bI5hlHtKgolBMlODM+9Dbc6vx3JOZY3eA+NlDuC
ieit7bvcm3P3pAotVIry5hFQB/a5vO2lyEar8drpbMsPVSgmba8YZ3dxOEolwIHR
rg5qhfVnp+urx+xax+/Bf+Vd30YQkv8CrjgaNN773P2YPVov1WgWyg3pUf0wbWOk
Z6rjBiN6rFsTKnbBEU1z537pacWRy8Az+s9NU8unF94litX6z5G6smLEzribnIw6
P7a/68A7jC350Q0dfqX1td7qj13JEnk44VUhM5CoXmwf4D/3krxl+FT6nRkdiGgm
T2/qeZ+m0IpWzKAbXG6biNLlaSfJuyb4uBzlc4qPyQteq1siiTEi48Pgn79Czqh8
7srw2APn4Un0mMQkcMUug9GQsnZnRQf8KrBPlz3OmzLjwILa2qEPQ4mUdlVvimyO
Qr1vVr2ziVnnEL168br3UUEQyP+5F1ETPguSxAEO3+MS+5IRQXC3VPIh1VZqMTMh
ReWg5y4Z8FeDtMa7ALuYjiqt3iQ5DkJn4oWgr8NYSFqirzgP5VOwxPkffsZMA7pI
zKxqHNDZGIWuebyEwkBTyIGgx3TobIiHx2kdOG7iz3p2B0pjQMjT9gcX+YlxPBzl
cs79/YBQXZzjXnkT6W8lFGXUECwRB6I0sw0wti7EqMP3BaddRsQ8hdcewInAO/bL
tN3beXeyw9TzBITkWJIkR8yXRCrO/smQlolgAKVU1ha+uc+oRSXA3P6ovDKLfak+
f9kk4JyPXKOUH2+t9crMVH27q/3Vo352z//VeS6NlCkF4pinz7XUDCgG7xhy6J1m
3Y8T0W15Bh+E5HLWvxklZL/+hTzCK5tIPSV8flMSL+dsjB5u/todd2PqF30pCANX
UYP8Kez746VLZRuZW8rUa0PR+df210OLbZYBMeBdh5Yb9EQjVficdtI4LvjjXhjd
Vm0dOdsyOPcoVNNJU3MVv5M9PXD4B/yMc/pOJ/w7ff7tpQ9WxTWiFD8DkcDm6Efu
21HtamDduUyaBWauqbS+bEO5WOwQ/ilH0P//1W9ryDdLkufalFCktmUl2Vei48VA
sZ7bSD40b61jUnTYsbS578Jijuwr+t/SntEvoBz4osc+TJgJq4ls85oP5xchbJHz
FAZY2tPBdjzo45nqniwXgXRgaJvFgWCmi3DRikLp3e+htLuL+sA97ZzntYj5uDKw
wpnh47fJMUXv6HH/mOR3X/l16pmnS/fd3xuR/257j96364y5+B08d8gLEDiDvlMS
suVWQY01fmFza87FRWgY6k6ITxk1YOokvDN9nn96jepLZ9k4Fis1W8HmxtngRGkq
4RdAeDcEp50ygskLAWCfFvxJ324QxSnXr4L/RlBieJBXYxwBZjw2/RGzCG8hkbjX
4y7IHKKqt/4huy2Y1518wQOb1iItRjQosgGVJYYpOuxcbGSTUh6HX7ogL5x3deQZ
SzYQ7m0i0txHyWgu5L/xBThP/9x9CVTsS7N0iCKGWlCHsYJDtQNA/tTONPYLAm85
1Hn8xfmCjzXfhvgZJGxrZhBkjp0bfmiAjJMDVBNwGOrf6UnryDZM9j7rn578vBD1
I1jeXMtzGF62L9D0XWeHscDOmL8HnJwGEGlFr8BcQCkkKU6IpJ+08qXtK5dgWJDz
sB8MQEwjZZTYmBxW4WHrhsciX8G6r4V+9vSD7hbIjboWpPUE/gzzMSjCJScf3zRA
k6a8pD0kXgmQvO+lFJPAClg3FKXuoTptqVCr8bFIp9hwlJQLh5R2g8AZxceF0pZL
e7GUafYf91mOPX14jg7sdkQiioFPxNKdeAfgbPYQroLeMDIPQo7Yfa4dPMvlL3Lf
i8YHRgeJpNsN8vU1jAWGNU1Ay8L+iqiAI3X4PhHPrJZQHflUWlsdi1cxC0xGyFSz
wcIj9P2HsCoNfc3jCUeCPQW8E9N3cS9ILt1WWIyg16QktZMxM4Kkx+vA2V5OYX2o
ZRzzWL13B8xXAJrURApijae0LufkMIYVSD0NQ8h+Cqr/XvtQpaqELZOMaRMcZKm3
WTlcuXo0PNz9NZoUPIz45i7hyW+3vsS2COiN5yNg5f9ikfxszcCl7xz9cNxvYDD4
ZDQybu9DKNOaCNEMIJ+pwFEufWG+DdeiNJxWkhCw2XeBmsP+En2Gp8/J0sUB7A0S
I7po1pzZeYLOUNK/m/fnuUugKBuGacCFgebMAH5ApEPgt0Gn3itI5SyrB+27Aanw
E19U3sQwRkcBUXLH0kuODKdIQQ5cpO4Lsi+Tw59mHVN8iOvc1b+qFDqG4kR0Ncz3
WqbPRKs6QCc1C088E8LfBE2y2n7J4q23AC4JRoYxrD1bGYJiS4Saq77e1pTEFFhA
c0x1j60Q/05YG4ha1zTy1NYuhRp8j+oYpnWnu0tK7cUqAFGGvqeRxyQViF5nWFIW
co/tui7LrYTMqSrNVRC0fG1PPUbdPCXXZ8KSHLdRuN5nCS7akkWZ5OsQftArudYo
x41wBUlOSbNaPlGYegkUoheTKtSJeJrMpl0MpXyX9zATLkhccYH6ftEAHCCzYnfH
WPajRPtDA+gRCI8WigOfXAQAFMV+jrDzBN95n99nwk7WXCaNJJ4sn6WXKLvkW2An
V+XH99JF2ZZ2aBY8EtogV7wJL031RrEVqutojG05bY/dnyWM/u4dDARTt2j6/XyH
LHTmEEbTQYU22VCc1bUuHGQaJJulYAULSllLM1pntrwLP0H43Fm0y1lWCTVtlt9c
zBT/IGCoIohrE1m7sT+s9+El4m6NDBF+Stt9/rME5RfXVXpdtydmkIzdW7SFH62o
g6wbSLV5OG9eQr43uJ6L5d8gWe42ZPbQJpEtK+fUEQurTqKcotR5wWNM8SAbsqkr
zvtpKpyZl4kIRSiMuK3x0nNVGl2PcSR7M4jhIXK8XMPeX56q0Vsagy9hPtdhWf06
T6Yj/NyGVpP4J7KPY5Z19dlVrPYTQBu8j/r1WMRIyYwoqAMqo/ISBm2EWJUqklzL
zu+m9Gro82SX7BUM7Xp1ePQw6WQqapTTaStUfeHhEs9418Dvwk6FhQX1oIRpTzxP
1wdNahjbmttlDt2nEYlXq1V+vFsP2tHmBW2Vli1PhASNT0N99EdJlhXBmBJez9RK
zbWF9e6Kbvn+Rv5ecHE3tCs8VQDVMMPM1VtnPtMt6zM7P/Nfn7E8C5EHFZAk1K/n
HDxMWdovMW7wprLlZdcA0jq002jZaCVb0mN09eK/hh9fOj6ue9d79g3cyW4LmNzG
okAWMA0um2Y/IHSNhL2hZXIu6AJSpF5pJr7LD43OvgzAoH+4JcjadB6qM2SANzUu
6ZqQznUQ2GxilkonQdhVm8jHKP6/4FjnrPjbjUcgWrwyUc7XqyZAMs7+rpYbzLKG
0yhI8609Za9jFyJ4ItAWX0vOS+xlRczGgqca27wW3hImTodvWC4c9TYwPnoeCKaN
cQJPmExjBYwVg6HzDmHBuEcg2GefDpTp0RL8Zoeb7sEDK5+v2zS4/ipGvLw7T7gk
um0mCawoGixgkmt6x25my8Xhe1X1fFxoHZYqecdYyRkhUgcQ+E4VNjEL1BrlZ1A8
8G/Njw6gGHPlKmyZ6ZGV7Bj2iK9IdlcmSsDy1z20fNybsR42jh8FzE32nqUJm+Ag
7G/Msiv0TYVI6Yvk5dFUJVBoWQoDf3DsU8/CR39qNBbepU1ADSkCCoeeld9frq83
P3RQormE+Iw8lSpU5Wwrs5+055G6Id/fDrAeQtYUGDSlHWRXYmBE4Ya5W+7sAI+q
R87chvg3v0ao7Yfq5jqpy8hTSOvrV5bPcuLVU2x1SUy2wzjKBiXg+D+IUcPxsn9p
1h/GZkq8q5EkFjsHYAfMZ1YYp3dKrsmwKVI7NYcxl0MuE9qLnWCEy12brJzFf/s+
ejDQmdG0lQzU67LbxCxu8dtfCdw8ExOV19noVS+zltFPYjJn6yp5EC1KyPwTY3xv
b2DMEavhxSRyJt2WAYepGLnnk0RipJPMN9MG0NF8V2mxSBXlt1LeUb581sLQHRTQ
wgsXrWba8NUI/lisLHmGUcJhTo3mL1J9woea/PSmVA2fOuYFLVwNecr1rHtSC1MG
BtW/J40aK0u9vtxrwoHb/lsUsiBjXkM/RfKCzgBKyYNQk2/tJgaVskrWYGA85kLO
D3EJeNvh3jK+WB5UTwNMMXHPw206GCVglqPcqnYxZV/VY09NtXr8d+MlzDM49vmw
MHs/aLzRD6YCD0Y1M3i3OyLB0WWmRCuYVP/55kleDXFHgYC+v66ew+1j9eA7Si4M
GMTvO/O3d+Ro+h0jycVRYGhEfEqf6PRwmMmKWLJmaDi5+ugDouwv2Sq3al2T9o6C
LRZ/At4eQAFKiXoYsI5o9BREa26uCDHMGk7ngZCkJL1JFkerEFxZ26T5yw71f305
J14JsbTDt7BLL76LFPnYDGCR2XEzvhLv1atWeG4YmZvFJ6lv+qGVG4snWL2wrcma
efk/8qBYHE2usDPUcJtPC/KyVXPCfvxcyyu2Rk2RNMfQ41AeZ0Xp2EromAkGnecB
T4js/RLK06b3ONcT9yLeLqS7NTc7FjTmNbpJaEGxmV0ijfdoF+p6guYpfyfL3zhv
7uWqqgcqOED3WhKBJYS/nVJAvtWMzcZe7qyAbDDtgEB43ucN+pC3ozvW8Tr/k0vX
J0fyw2gShTnB8BILwU3c8RbAcNZ5yAQyL1PJfHKvZvln8iuCxmcP/k+FXJB+rjBI
8rkjrlFhG2kttzeq7T9kqBWzuk5znu/FYfDxLF3vDJqp1yGj8y6p/7IE9bIBQQO3
lyd0e1y0smIrgfHoJ2mZk1HFaiTWpzk//OOe2EzhvdAtT470O2Gl7MkrKCMDsQaL
HhB490h3QPpjkiJd3WjG5VBKaY432YzkSjJprO4rMRpfYFnWZV7EqiQO4RGg4NfE
jlw0xCt9h81kCcZCMDq1OuMZzvle7yS2yfHIXn+ni3y9CXh3pallYIzl63c+5RQ6
u+G2PwgP9vY7ssM2ukBrlK8ZukiHw0Yj9YswPAjn+CRJTTSPIJJUUKjBOpY0pKBw
XlqHCod9gM3n+7N6TQfDYsLz4rGW9ykt5htJewhsMPtqShhyzx3Wf92W+H5tX1aQ
cDGzoj2MytkL2hRGW8HxUDvAq24zsu2c1+w0U82C8KZKltlS8vMs6/clogjJGWKw
qkpxn4kwkz7eITIj4ifbuWDJ51Af/ZElwhU4Fu0c3sr7J5qOOmoIpVd+jFGtmWaW
8xt1fTNPRkCczeT5tFTvQ1c3rkfC9jrgvDyKb/3MdRbTmdms1VAU/sYYo5pL8Waz
1latqwz9/cS95PdwnyiyJB6nrIzcv0XzU1WO8GMZrswP1MuFwGCEan5Fq/uobxST
nSywbTSb2CWdzVDoJ4+E73PDAV/eqFlPqhYl6biUAljIuXyEl+WbPp14RMJdXBcP
R597G3ixYH6Ds4vmUaiUcbhMa1wfqnx+rPU7jDJdhfof84uY/mERWwvkaM7Vhi//
fkXC3gf//YwXPdOP5uCHuYPjFalF3R0uYlbzQZGdWF8Zo3wPiZo8/dWbV/Ywuj2z
qt0bSBn0LTuEfjYjfmFAhk7Xl72KFpoYOh4+GEotatGqgc0x04RK23A3b5lWNRz/
LecdwzmpQd1vyIqim+Hk6dUFHFpn3e7iYAk8GmdwUEDWNnN0x3mzshKnbLxo07CK
G3Gast2FHt7kx250vAFtGAXwz+K8FZ9cyleJroUkQhSmDv6KxmjeoWZ+mH/Ttl1X
Te7XkDqn0eg17MvihcTX4HwNIrVnGXk0De05pAZPhdlyc4/lQCVlSKg5dioi8Iu5
5QxNn00nWAvsuPOS6eWUjuMu7IVSXf+rJXGL+k9FcK90nNMK3ro4pfHRG+hZ+kSi
T2NfcfiGs+jY1ChG/FSAjTySx7IGI/33eBlKxJEnLU3aE3QAElpFVfCIcnYocFyb
gF6okXSxXel70bCxVEbN9GqfWwifWN8vPF/FgYF7hI1nxoTJC8qCSedXxQh2IsDw
BrY7ffmJdGV0xJnFYZ4T5vfafdn/fweU0LYHjSgJEZ3Sen9hF7UYtAotnzoXGLIj
9wOqvUwpB0bnC9KlXncwiJCAPf756l3IdJrJ66D4hrlW8soD2udpFvdxnfsJos9Z
EMHaHMfks6uoOTq0wwoAaB/q0vSQJUCsMZarWYelb5TnMXyFk5UMXfQDDnnwRKVe
3BEMMlsUSZSq+gzB86WHVapqrzZ0BTbCQ/KNusX9dxHtleAlLe4wRGlMbqBPX7kx
Znck4DjxGzlF+zsRL6o8Gc/aRsTbE+PJ2D5RW1Pou5bfySB5q7ZEdMCED0HxPqTJ
26YMwZZ7f8JshKvVLVOiuF7ttS+sEMoM8ZFk4EVSX60oO0RjsmJTXUpOkDdZax9M
aApcDFP0P/66bhqOQpo3mUAVhRGds+p3Ssai8JV0rnAzs6/J0dDJhkuj2GNrP5PN
iBhmqIlRTHSfnrovHsBZVI54Hj5N8B3JlTqdtKgTfkLhMn0oQRiMaXLtzS7rQWsN
xg/4GccalbyljoWa7poLyxFS1PqV/CwKUweMp9jBsCZmDkNtGOoA3Dy2ykl8Qdxm
uv1vkfJBsCd4yFeVJcUUjxvN0lsfF/5zDieiwB85wQYNborQb45cBQ6BTSp9qJAi
lHNwR8P3Ln8G59+A8n2QwOX4FNhDHRgobpeI/6moZ4zcIYueEXFBs48QIkz71YWJ
44ZlOquDH076Q+5232GHazy8tewZl+iIy8CMw25gE17sNhFUBzx9HUzyftLQiixA
3e64d3GS6lPaUa0xwcELTkGJ3iPpuyRLsg1FS2XaanOTUkzTPfqHtHzvKZAd4TH8
kX6bQQYs7f/8Yrx8k/NP7v5iTJCELlzGOzNfjNvu31f8jo3K9aYKyt9m6pk1VDJE
LU5fb8wQnOPmyp8PdJF3++dKRmjwFDMc7RG3OGZ01q47aApsoyzpbrpmrBNG3HAz
RzahhqAMx3aluL6rsGejkR1mVwyRNWfeB3RbMF1tTZJAgAnV4zGzGQlosfItrxUs
TluP+NKphQw8ksMMKMX7AIOpR47KDUwF4t6uL89yg1hGV2uwo7KzkuYb01ObSOJJ
VuK+RCol69/F7qpaO+n2+9YOJMS7ROmu1kGfuHFMQjJK9AOu1vBie4j/ZQFMytUc
sJ3iiZzsksyEYRUkGkOkKbNmxfK9DFVi2n0Vhg+7Xyis2Z3j8g/ljg9h/iItiCGk
HAOPYzOJG9q5VRxhXmY6mkqGSd+8JVMNv/dFTjPnnOag5m4TkPH9iTrrrH4Cckq3
xFsR+Jfol9N7b1t0BwCJNy2X6vsrti80Sn1xvN16FuuWVAAIEPJIJmCGhkEqAEiT
IV2ptFQmzYLeVwcK083p2XXPctpwWEJl/Fh60ym2NUnQVO8HPHXha8TunS0zNC0h
ApHbhuSprTBpkzCCjieW/60lyW1Luga5o86yBS+PdRL9bzoAWJfTiFA9F9Pp/sIr
t6ja5Pf8qogrUqYVriY6tjLnImDvpHLMgpMX4eLnGITdQsMujBQeuKb8jU5NOIcH
MwBgP+SIm004YZEYaTvCa+rQ5gzuQzoFHLZEyQCu/x36X14KoyBezocPWXURWS+l
eyhJxxUQ6QCIT6vQOYGfe7rKEOTlWE/zuibLOm7U1snTNjj5gxUHkbmzJM35JkFy
9JRyq2u91Iv1IC77ni4iVchDRo4ZDRuIdbbbp/FveQXr4kL+6PyHbuxanVr/vQDj
4l23YfTbD2Vp0AAlIGNqo67bfCzJdCwYQxt8NSci+2jXKQgk9T2LpSpSXnTY6onB
NWplVsuqxs7exrzd/+cJHPasSY0IWb7RnbUUri7IqpxYZCiT1MI+RrtyKXIkbfWn
zjQp326nTsgYZt+RgDC+zTfIiKHIkWUr39FbzWzNYMWdVjBSKrcl4Q8PlFJooepY
hyY8Cdlekl+oLmOdSueRr4XWOY76WiKenC4DY/v+wVKJwPoDtA9tDyw1VvNoE0MP
NvPs+z8bN8/ovO0k95LwLrl7O1lwk17UCv2u6TEZbw1RKwa3BaaheuysFImGBeow
InsC59tZ+7GeSHg+McCEXVi5mmlybFahJT7Uci8Ha1pGeZlHItjJtFDnXCfdxUkv
xICE1GcTWpVe+cwHw5dMv7w3PlPJGodNwac0kRDPQbTeNKFBaSo3XgmR+/YSZ0Om
7uTHzw9HlN0buftq3azKeGI4cAKBIFg0bKUKwWDRyqT4ZURdLW4rKsyVPAH29tcL
h2vXvLVD97DGm/vgYIp7dz9FuL6COHfW//4aEFflmFXH0fwmIdgkNoLqGo1c/Mjl
Mum+gT+R2mKm/Xdn5HnTajVTCrw1Qqk5If/eWh+DNoF/4ComOOu6jAFMdCE0Gk/G
hGlEGJddu7Bg3KiYH42LYLYTCf/oQgA2WorHulZv5TsYdJqdAePRUFcFf5ptWHs4
/5Yos84m6/h22Py9i20Ghhu/RQm3oUPKAyVmikXYngu8Il/sfqXcmQmecedJu3ly
JPxMiqhtKf4f0TNkV3cp/hnNSWquMPn/Yo3CK1Pjg0Xf5OySLPCr8U/nNP3PPlhR
JrCDpQKUs42ESUSoxku3qY0L7djX3tpIinU3DkrFUnkjQsb48AtbTeWzBNvK2nd7
PXWGmVyJhNxnjB1PSEwwUaM07EKCYZEKsr4rcVH/fT3hvSFHAS5gnmV83WEoggUD
Rqhl2qIs8r/4Md2C99GAHP3XP7F5/tOGP/QKF14EV2dUZTJT2IRrCPeSGy+YKHox
hr/sfjq2PcN1QuVX/zyJwatdz0/z/50WnxIvc5Ff3VLxx0xXdo9XSlfWtFaVqrpq
1h9pTCegmzDmuAJkwrSwz0ptkrKzKmNCkBkKwjmzPiycUi4iCoE4tGP2vjEJt/Xd
9M0HqwleuD2IZUEXHR3jDDd+ZFVXlim8K9N7gbwtwPcRLsDN/ERLiZ4nQQetizM5
QopEDcte/Fdq3wQyJ7E3hFm15NRMaUoVGWr9PrCDEo40M2Ntz9Vhwjy7zwkfuoqy
fKf0kY8sQmjaIOm9CvwmNDNJXXqY+ncEfKvJvaql9sZpGZr9FGxDXfTmoJ14eP52
sTdaA7CL5nk6hclseb56XxBUvpV8Mz/6Yqlb3KF/h09vclbx4nQpWBoNr6xL7/zK
JJLBoUbzrcBgxcHqZAHt03MF8Czit4TMDRU2ABHXas2GDJ1v+pWuDmguL0oT6MIQ
YN1oKbndlLmxgZzBH8e8fCwAOZMfseoaFIQYLxGrf63eUQ4wNEwOzdx+Z9cIMwsq
qC1BD6c119cYJigc+1tbsglrxLxF7GRpNs0FZXMBdRnaREcBMYPl7AuVHHYgo+aZ
SMTvh/SLbYPjLoOCaGsVx1CSvZEbJtmlpvrSEQ0zV2z05RnS8LqJPGAkkxkhJEFk
uTm88KkpX0ilnDpXx8ijCaAIr1VtuaFGNRjGrWSvaQZyVIUDLwosLge4gjwHOyu6
wUNGRbndpCk/Utw7Rv63XRcprUselicdObplBOVZog6GmJuputVujkVDUu7z1IVf
RHM0HDZcVEutcLdciV+e6itn6Dt0i4l7TWJDZnHsGGGVvt6x2zEPWM03D+nkfBhB
RI9snURXj0LBobUaWNpFM9iHeZQrvcQFxHPxdnRWOfdeOKOzMnwT9MAcxwup473H
z35PZ9GKBNmNtttlDLHfcD6cElHloWReK4LXTnibOH/nx7EDd2H54fOUJqoHxXPz
BTsWAPcR7+giwVjPTDXS+J0aU3aIdztIXJzCT5KUZD3WHGxbETOieSey8yF+DFSy
zyuZdAXSeI3dmhhELF/4dnEWcYxpxkWsjiJn87fNtG6WLWWYNw/z8ZNRepC+3SHv
VSWjGxsvLMecX1v0MBP77TFvr2nWIJNABXpuexaru5MNV04pACZa+nVbJVLbyfUi
LJXph7VrytP4rU1p48qMgsGYV7Qj4neAmCXV2fMz8dK/hJkulwAraO9pvqC6VUBx
Tx5kPc6Mt14WS0CWY2awhxZ8yPOyycR7B7VukGlEvQipeWs4g0Xi4zHZ2jH2wS6E
Pi2W68KqAusTqedT7q9EuT/4/ll2OBSuI7L3DG/XRngif5lqnJrrs0d5m0rM51c4
A++6E/9jcz1hJ5nRP+FtXtSZTGJYUWIKBLNVTp4NxADirIsWZazfCQMUxCKVi0Ke
not8iAEk1te87LQSUoHa3H68/0btz86J75Mupz0Vya4Jn2k0UoEtVqAREPLlWJBf
beR95DWKnqBuSSkd+WPyGy63ecI11G0xQyf1TViYtcDv7YOQ2MMmyAV46bpPgjmR
HgxEneQIqmNGV46dKcKdYl1kOX+OU5GCntq2c22tw0ghmGfABRbhrH2uxU64lw1G
ZVnfOJPrmMtu7ypJEjWWsGjbeaK6lTTRg9Uu7tZ9pAZfZFMswuf65xlKhb/Pygci
s97/1w55gu+vL7PQkn8fUCPvCbAhPj+3B8eQn2M+HQrwkBov+VvdmgebrZuVYrjH
ft6nd4s4TmdWmD6yMq4OUnpCcVDYNZY5KM0wUfFCbzugtc4av9JF6z18VF4rMhpN
oSADFDJxMiUiFgWzJDP1zaLhHFzHck4/ICkKR18Dr4BhH1yqFq9l7byKGI1ARiJi
KHOHjRRJrBfAG7p2m6WzcfzayPfv6wvGW/77W9Y38u+aSAtlIdfWD6GkXmSJivGC
3rme2MzmGFOrpDsoQoVjt7P1FUv11zzHK6IbOSIexcucUCcAHI/nuvaY2Qp/AKQQ
cgeV840y5T4FTpjorMhd7+qbsLL3XnwHnxG//D4lJtW9kIaZwdbu7awaUdxf5Ol0
IsgmCk14w6AYOOSaGzJuK6r967k0JFeGpdcWp2NOoKUoseJMi1BSodcwLjHf8VrH
6kV/M4WSsNBxbZxaLGIUWItjO4crfijoP2M6YRgTapvMQGfxDci8Ap6xBOwK7YKU
zypzRv7snvgcqEsJ87HqdR5DkGdIdPfLY+sHUYhk+7u9ofcYOcDgaurHGTJAnqHf
1eF29C3Dv/M3L1md3lbIfY+bFG0KJld6NU4CN56P8hsAj5wV8QNxZpkLuiKzZ0+f
XfZ0kPXRym+Ce8lfMIJ3Ko+gfzhZD76JKuCU2nG64u9yiXW761jA0xUFQwFwj840
ZekkYgSp2symmuSTmPC8u4CqGZQiHNO8moVYtf7malhXw55UUHDcWECW9EKkWvng
fVJHJWezlKJVBovd6aiJ/O0s3d0GXYfedmOT1BRGDM9GPJDTO4k2AfyO34z+o2kn
LWVFvuG0knVnWlZ6tGbaVfJgTR79hwPv/1bKKfppAMxGhqVWHkqLYBy/USBYeUmz
oHdPdqldWvOvUG/jCjCAg9dmbSz09kCgaIBewYlcUzdinJOVkM4An2Bgv6wgRs0W
7cls4Y/PG8mtMOtWJC84COVdExHVwSMbKu3Xk2R4QbPT+2R73oPJl3DWCpTO6PcG
/WVmJ65wgkefm6/Yx6onWF1iOlFPVb96BItquJEac68XLqAYsT+kpoNHQ5Z9T1Z/
KgjtFGRw9xKyS+ybD7oJO6THvh2nWh0L6kQGj+UzpAGus7V1aVsjw+JxpOSm3n2h
+YCIQNS9+OAxslBUYwIzHbwv4rfxIFLpdq4P/+3ExuRi9JfrLotj6PSXV5avVq/o
Mh/uDCx2kC5YvYDYGgukxYuzuy0kqyIohiO4popkZjZYkLJ4p+JikxZ0M7/zse/o
Zo7GpgS8n/IGSRBl4q5YQbuHAmPpDigpEtBSHLNmVqYaZI0HJmlYBCMt3RvVk1fw
8rptbnk1+mFg7xR44kbdAnYN6W5WClxgY7UDZiTs3R86M7TsGN3JoaoedjBJYQeB
MVS8XxFFfX8JzXlBGU56ENOQistReHar8r84jlneyr9iNgxfQ4iB/cmt8PE7Ckwd
YHnM2FrFLOgTT9TdhntlBB88hUQcYJCtx1WZEvCE+Pt/iAgAFGuSMMNppurz92eC
BWtX8lFV9cAi4u9DfDsu0bg7U2ALfLl0R1zDyPUEkB1Th1E9cj6wSlZYTWAxeBWC
h6I3CwQdUN5NWR7aCqTEFpRd5f3aHDvICDPmPek4YYrrpiYFGpk4n43UsmqBkkhS
g6THYSgz6yY2D5LxY+m4TymKbVbvF+zyHBs8FtWJLZCppnzK6vemiMk8rMR49QbX
uLFzpTcjOX6gF6EXbMSLDRd+YPCDzZXt7jLKO4aopBClaoY3CTLFq/TLT9C3YXjf
aBvf9c0iwW8vCpLb732hAaQsNMmKH4SZSNGOvph3qvGCQfEyBmF2NjdaJlJaUV4H
8GJfH0E2Gw7Gikj3sYU9WUSd1Xbi0QvGNRP2BS24Ce4re1gZ3nvttNdrvUfe7Wf/
EGDFpJcW7614Gm3W0RKD2601c81RFKuRR6dTX2g04YKW2SWi+byLGjgiRHv4D6P5
Wqv/+2smNq5GWg+Rv2Ehg2zQ7lw5Y1OdPnXrb092kCwLe22UIPxBBx8sF/qArMR3
BzM8lAwl8q+M5oV6R5TlX/zG62tZw0dHifnMW8A6yEBGnrjDs5nLUmGlgPprTFKv
KdnMCYFSrJ6LpZqmoO0A4mtznbslpIb4GBU1eP7yt41w1E9tta2Tldcg6vFMsNuu
D0ZXYL73oLVbP6b6324JrdIrs9WPVbmlbLd3PLCMUc8IiBlr1pHBnI3Vw8ORdZOu
TwtVMG9tdi6rHAbUN41zI+rfkxMKuXA1L5wCBZX25Dif9La4V4uKr0LzD/gU/ZK5
W4rcq0dPKQNA61/fnHOHf2Y5vxgsK53EE9kDYSfiMKTUOzWMswAH8PicVSMTxvi2
3vnBuAMTFKOL3Ch9KvAw/QVzozxQeRkQrE00jBLWt9R+H6eSMAZ3dL3jcf1skCqf
5C98colGoec866BsflTcIDZ4TCARIe1d+wlPP+6v7uIDvOx3KpZ/tdY+2O9OzF7L
C22vjhmMlMMJQgA8EC9UYpMfy4dwICM5BQxe4Ry1COVB3AIF3QDN6hUdww8DE5YO
fy6ZhPGCrg73ehPIBMW5zEk2/trxqVlBCwvkNiefuj2LEyrxyYLduimjO4kQWBh6
JTvSLfP2Uh9tR0bKZrPRkUpBG+6N2IpIUTvwg1zT3EFTt+uDvWdAck+x6KGUBoMt
M2wqmEwCNR+fcFr6o237rdYUJOyzsipZ3unpZwHP/+m7neAWUKjjn5NBYXwXCfLB
bo2a36wmlIGyUjMjWJTqCWOKfpjrre5sn6wKn8CU5vHyTlh386oZO76eJFuMRo0X
ff7VZOD03MWwQzUz25SYSzhUvcw1cCGg7iHTuOPmRFzUxdZGEH4fGZUwpWB6BoVp
5PMwUBYFc7ebXXR5aANBzhfU4bnW085y/08/v5bI+0zdLWVOBObKZGGkr8wPk/YE
Dj2Q/mQ7mWIuhCQrBRw7jytgxmkDSoufoGyvZR9mgcVdBzvPnFTfiGWH0wc1J5ut
OiNr+a24td0WWoUHlP9o+/CIVOoMXffXVdMh0+S/Axg3I5VK1BZ5JcjaYC2frqZ9
JBFyVFC3/M6GZMKqZQHUa1/o+jB0PmODc+8KoyQL0/ufD4gdodw7KA2ep7LG4uAq
UfVGMRj7dY8lFx4lYP7MigULvrBOy0wOV9GtmscU2WN9xbsyEv1E1oUYqPCl91Td
U8kJGNHu7yBYpIZDwhLQinSF46w3Yk8ktakh9JcCstuSDSjwSRTsJ2Al7t/RCX4P
+EuNFUR6n8Bfoyn2Rkn3MmB+pfKTHiVQENt/bccfrl2myrKxev6WhFf8eBB8HGoQ
WNzCC1CCprCnXE1dMOLnPHVICRK1uXH1dfFEZ8DDgG+NeKQPln9Zp5Oh2YOS2fM0
nGuRMq9nVc3XLxtmiwtCxLLKGSU6huglGriU1i6JjqiYf/oiWM5fj2Y5vlibpFTf
k3g8bYpO7GRfIMtnAYcfht5GmLA4ARiWjN7SGWwo7SoVNINis2c5ws7bADMdya5A
hlxQQdkhE9CCdNZYT+LgcljqUgu3HdrQmGeKvwEM92Mdk76iBn5cpAMtwSljZ/V7
dP0WXuSV4CXG6Y8bLp490djnLORczZ1IWBZ+ltvXFaLDwJoicTVLuDjb61kDuS1a
UfbCAFAnYwfG3P6+cQsckMR7Lx9fvcjFt7gh0p2VVv5FuuMmJ7j3lDgF6F3rTFMt
OMYHGb2E1XVqCxxAM/m9Bx0X1IeIGBNaQR+ZIg7rvvb9t623xCsGVNqDg87TwhQw
pIeUzS7cWF24iKQ0SGkQkZ5qweiWtpLiz4w6vfl2hRjWRcQ4MHO2XCux7r7BZWYh
zGTHMTJfFPGeIjQD4f19kbd9RThyKJTY8o/QGkxFCU5aMhlh+XEs+gvzGCh/1y8Z
7T5tGRcfbWeOhgARzLXUwdMJ3a6wTPd9+xrpuajOsEr670DuwRnQ/Niy1RAuWu/Z
N25TTjkcFTdTixjIKRDQCshw7q+Y31KDQomoj5OxnsTZ8JkSqy83Qqy0nz6QqpDK
roXFWkHl6nNSD3CcbGUluDOxFeA1j15xFmw3q1oGnj5f4tWGcjS8H4lAD3iTqvfN
K1rgbAxnUyLXHuRJzvt/Tn5tTi0dW60M/8euG5wmJSQ0VVWe1AmbUpmkN1fEEzIL
PI2ETOeX1iPOPWMPKNuxYn+iPJEACtz86TRwp6hxku6zGNEBSILWMm4ifZ8MLwY0
s9ZvkiyyVKp/vNky56Gwv4lcFmB5//0FcybI+RI6S34/4JrSpJBQ04KV4csyp/+q
LvAQ5bkfVgjneW3vbr4+FDkA1Uiw5C/1JQVo6q8Yl9ERbE6FMutqwVqZvLWIIfNv
z72yNedKAJO9Zf1fEC0oMf/wa9eCuu9dUlvBG05quAzEMZrFgYY5PoCgz2MMeQ3n
UMOAaPh3ybELNRLEVzPDCXYygBxJzjPesY8vxCP359G/kUuGl14xOgycKvNktbvV
w5xASIqlPXtq+dmXnvnCalHiq6CTaUlPgMA5kpTz5fZHDXFSOe7KhpyJL961ubvn
p39to0S/iEe/+go5IEutDXtlOTlOtovAPr+x0k24WbuhRXSdgkyNTGTNX1eQg9YO
YiSwh+54MJH2WZWgmc3gqJwtoVdanIU8Yq7fWuPXz7ul+14HAokoawJI2JEDSF99
tciCj+Ay3DgEx398L7AwR7Zcxbnp42JU5I52Gven4z27MPr947Wy0SNubBwDwoEV
ugICShlkebqQdJ8hEqs/s0BolUKhrvY8dB9lc/4BQr7AyZKT/8XFASJRqIZ0cnB6
88yQmF8I+yf05x+9k82OQlnTCnbsNa9kFXqhcq0Mc/R1jVfw8hVUiwtn8FsKD2N/
02qklDtX/1yAdX92P31mJylTtOHGVuIjJMQQFI7JXXVTVrHLCapYiVuEba2cjcR6
aH3cVwHUjXd+oP7It/Fdau0uT8S51+8JD8TgC13J4AtGGzV+LpsKz3a9o5FOAJxL
hlK9SYwo0tH0+tbonZMPYaYtZA/4B+tgIbF3oyzFSx80IfQhhgP3ijxqkjlaN8Ld
e+pKykXJK19cYvPW6nQe7+0NenqWv7RnwCea+RzvY1B0Sa/J9CI1X9V2wdtoENGU
RO6e4UeetGlY3HGOj6fq6pOKmoVcg0FIr0qWCE2jdfAf9H5wLI0onvGwGVMo7TA1
/znxjwBX2cJ9LbYehujgVwtSLzom3wlVntHXPzYY+X43Xy+3/Djtg4XDp+pMuga1
wyPr+tesrPMwLuoub/E5woyR3kHqVhK2+YVuYLxobcWDo8w1rXmN5bHo3RZbmN4C
blxGCWjn0BB2SIyn6u1Hnv3T1lowSK7/aCPYBekCpi3/8HYKNOdYJMSVjRW0ekL/
oQ8ZqLFQMt9SWg2zCaB+96YXo1yPq1UQkUazV+vtsGLOIlt0fc66qPCbqIqi0aDT
5P4mlDBiAjZk8Vt46zAF4wcmpdw9zhV9+T4gOptVlTMaJujy4PtnltRgC1jz+cDu
QTD9oZ8eSipMCw4QMDMGAQCccWWS8djUq0JBrP8XzNWJ7Tu27cKqqirPJgNnWMIP
+9m7vIUnO1UM9xmzcwTbgPafx1yCWf/3MvO7EKOO6hN4emLZ8C7Uytbv6gf8llGJ
1BthCWCvur/WSLo7hsvOe+JYUPQRncmOZSpaCw7fJGiLgtOFf5zAFdDUpRAsPon+
ATHZgm3UDfHseVUnNzO+cZHLofPh5IIgViHvw7/en8hVd0anLfiwo9aq03myQ5fS
xFsz4XeL3EpvoDfVbBBMIs5aEDo7mY1iP0nqgI7MbNOCKGj2gwFv4B5c97y9yU0T
yGePeEHUrkLQrcxJ+zpRBcdDsmcoPpdGsQFXEDLU3YiQHqWAxJDyzPmANPuKzHHT
bjKenKd4XXmJV8Kd7/BtERt/kwr4HlWt/1S0Ta3bcY7Zx3Y1kPxw/1VSpFjRSBbX
6p+l0arqEl43CWlPvCReNaZg4CtZSwrLP/5ej97NxAEketNQNXqIkMy1tdnQKAdX
uPH8hmh9c87TZk9I20BER2RizLpOQ+jANtrggSAhrIZNUEnvUrVBUl/GuJAnDpM9
HL77vfBQC1PqreO72846cYk5UyMolGVeB2MS2UVgNjh/dMb7jRQ1xJW8NHU3KByH
ajf0dHYFckeYpm1j2Je2g3y9FzlP2SpmAgiKe2D6UdJvk8naNbnIKigbDL3LAmsF
Rj/fkBUEqCr7iEPw4obGY7D/b87ei+q9OFNgsiq0JvWtffxhwMsU9xgKCkwzO3H5
ubVjuXRBVU6TN26udcZ5jFHrvzJQktyyIM6clWRA4EHMEx5YdIe5jKHblUHliWvu
z+jpBSIxvQv+V5HRbqXe1XX483Bh6ZzBABheFJFvAeDux8eakOyrxIkJLONkPfhC
ldwH2HxvIcE59afzhIPap+xNi/OAjoR9ZgpmMhblvnmasUQR9zll103+FTPERIvn
SK8g44nm/hlxDEJRty8uAdToUM03ABvng3cqpSfQqqViQ+6OtQkwaj41d9wmLTuj
aXQx4NlxsAitMnxLTB2kGpNlt8J2xW6blo2Vmld8ongONMOpIcLWnaR6ASGOPBrv
5nLSTkmJaxBfClGEozgWoO0MQk0Zr8uGRcN66j4Lv4LMuByyI9x0lb6Jkg77Je0+
tUHV+oiiKZnoc5HkrdPKKi/aKy0q5YB3p+CBL2db25DIdehnrzGm6YAp7aDjh2g7
aR1pGf6xX3LgIxHRUG/4MKAgR/ReT/l66KYaCMHdYktlj8Dl1Hkt0rzvccmhz+KC
lYX8w1f+6jn4LZrloKX+GRK74ku4fr3BQkPNfPe8tDacO3v2k5CviXzfoK8FXKXP
CbRk9UmhzT0zLsh27eiNMm0d8ncrfPXdTf1R+brjenlbxJiSipQs1Np3MIz5kSlY
abxiU4U+m3R0e+BZ3kMlGtwbgmbYL+yE/NkZMdQ+EFOHzDtsNMdUU9BxSAHnCibc
8o/UR4iO/pYq5XHp7taB2NdtVXNAD/WOwAlpmhVgOFvjwc7ZTTiIecpUbI+WKQQn
ZabpbFtNCmTWinlwW4aoyf6ko+PYu2Z9CWM4q6dv6gGJFrevv52TuoFAOr4eWnHO
mssFiePyCVbrUFE2oi7bfToijEOHbSisOkWWtL8P0KyPn3eqoWSyq4+2WtY11Pm+
gibMsie4fvlWY4ETNtLiyIaLsHq5o17vz5jUXgemU76jLRGZ+8yL8R6wS1MiEilJ
N/xNp6rjs2sDhi4L/zAf8QwRwa6MoEb9wMIPCLuV3N91yDFSM/IAzlcIB+iMiicC
b2773x/vDFaPho/4xHjYIiaCSgvIRb5cjgu0ag/iDolut9GsPtTz6XveCJg2hqO3
dH2+KHqYyK6VnZoIDZ8/w8urajIzsnMTn7pznmO+7WdBCjYF5T1UFp7uiFf3f0uw
vvqpir38qmOS1j/OxeYnRqoCpoT5QJGmKPxEm5MychJiRU26nxOmbOExyXmbCaD0
YPk4yIJyw+rI4+gdIts8ab0IUHTHA9oElXfq5c4kZulF59YjaAZ3fVdC9pHlxJiT
NBRd7MC/F0b77N8nrvJsbuk/eo9bhq/+lRSHNyjUqiHRJ6KlxnyLmeAIOkiEdMq6
HBFM93x6zal0DQEea0XI/dq+Ju0ovzxbuwRDIs6BI6XbbAJe/129kClqQZo2W46i
8W3yIaXGrh3wHXNIu/KWrNb051DNcpkJa1zcsd00Q7iT/5r70UGWBScL2oexM1ES
qwFC630u9rSlKaceingkC6/eVyn6K5f1KCa7om8CjYQhH6z5XSyFKLXRIsssDYwJ
lL7R/rPgFbsQ8kmjSermkF32H3nr9vJwJb947CpjvuGtO96OPKF4jHjy/V8CAKoT
35bysE4EbXI4Vj0c8vSJ5kRL4z3kENJL9HM7gx3vISRKG7Kdq3SsDBJWwC41akKU
g73g9mFb02HnHDEpMKw5YFREM1NGfhtXrW2BffYIbDXoS7vEF/6mwiGk1QWl5fis
F6RCoFYDRTtF4+4OI2rbmHSipMdPq07RJ2i7QCk7yKMoUKrDnAsXFL5n7CLy2l1k
jbGhJn6QM1OKuje4ghdvFNnib/MuazEHrBZFdnNhM8qLICxGSD+dqovn+QWo47t7
RNV9SdjykaPQAtoTOZ1upRXnpf8FcgYqZpVU1CqNUFUaWgJcKeN+KHZZIK4fN+j5
7ngmQ3gsld8XchIqIBtYNkPhdwYHoV20xt3533m0wc8pokNnIlz/m/paTDECdDzJ
UpD6wrBuMEEDlGFw9sBpZ5GLA/5v3HsCLW7z2DfuXBahPG9iPpfhXa9i851oSNN9
ezZ18Y3mxGWe1mypGNzKaOSTFmjAgehT+N05fpBUMQatX53tBCCqClaAvqleHjwp
e/B6vIFoQEQ9UGANtFEoOJ8U/IWaa1AsQOIsFKJwS3wmkYVH4HtWbh7xmpFIdbDL
/iYZeWLy0UDDT2vpTFOYZPgYRBUypIEvGten3+3OPfQejmq/Q1Oc4DrNOgBea10q
+F/1fK3wMcHEZLfkgz9JXRtDgjRVy3ZtBA/1HkqVlwpADH+uW9SGt5v4zQXx5DGT
/l9v6sCtvDySPUI6Lv0COOb2rT9tBWa/7fGTYoAbPElFUCgc8hxslil2XP/sanb9
VahS8wnPOcxHC7Q3t0ctqreP7x9x/98KA4zRvSa0B5lyWDEcTgz41nO6bJtxIFA7
lnMXHOcuu4SNaQQAasGee8MDly74CZA2tnbizGsXEraS2j2N5Z83cLGucBl1UEUd
ltwGXAUkHNDQE6/RnpjUX3WH2lMjYG7k32pMql/f3OJnUAaq4KN4cZswym2tV0wU
cuH7ffukAZ67HFlQXfmLcxrnVuHo/+O5VxAoFr42fjoa3O3PSx19hwedR1mnFsiS
yvR6Vp3/ImMTGT9Ry7zsyttftSJPQ5CqJ8v9KsRfxnMSO/9YvsHPKJpivswfb6T/
jMY73wa2ini5W2dIa2X7JdO3vvL2dIqg+wTtP4H28nHPWPAjvGLhbdnkApg/Zrj5
FpUjlD0OI3dz9k0mP9ipauWCUDPhVy/bCnKdyDD2KQYV8sKGb/MpL8nT/fPMbk/u
rIiDww/gtnPPWWtyPNG0vqzZHqOGZT9TwdQrRsparbae0CvkBYJj/GMpND7aOg1c
6M/fOOA8yembCqcd9Msu40AXkoZd2j0JMg2FqQowAwhBzcdDPeRWvh6YVq+AnVOs
fbeBHk9zQjXmSLdUF28+sy67VxpmO+ffr3p0357Fg4/7nGgZRHUH8PqkwATX9cuN
zxxzpAZkGDUxXwcMOwLJYGiciTSQJ25jq35xcw9ws8R1cFRaeOYay/dkrNX+iuHi
82vmwEuygrJ5LN52qE8J6+x1Ce5+1G57J9+o/vryXy+vO95csLPsgRHvoKwNpDaN
4AcTbKk+5rjMz8+suc7EU760B7G+AeoSEPkYyN+lBmvbVIv7CjJt4OLqbJ+yRxsY
CFYaX+mI0J+J89hLgpEqLAUXAk4bReFVpxsRQIElK+UX8mC33I+614x+LKPkqk3r
7d+AA3669YghhTULbkAqTs1UoOHtKSMafgVGL+hmfBL8XMvzmKP+XLj3BlVpp24v
IKi0PQvmlFSwTii4uF8Sz597ZByrrbqLnAfa0BaQzI2d+PBY2zkGAUz7dtmgdn3e
QnBdkH1cES1gF9TCQjTepIU3PCXOqfBlaCVxxc/HTlV+nui7gBx3RF3BZzSdpbDq
aqFvh2RcmqAf0iwUF1dFtq+HL+9fpG5K472LmcE4A7JwBrup1kj/0SHDEP4jI8tf
PVD3NxEbm87yudWP8gn3VSly+hDFEsUKHSbDZ3RTSSglPEiC1O8jvyFJJOkYi9GE
1GGWNQ+QvfBqH9PaLTcorVWgsZs9DYC1U8HB08U+/wST4ryOrzfnDZnF67vALL8F
U1roQZ6XZOKv+tAbd0k1wIsMhlIcDaQH9Tw7DN/Ncfopv4FWPZ2flh4sI+rjL1JM
oluAvl8MFQIDu0v6+zOYUeellnNDGxWCPB/xIGgb8vlYz93KVN0zxSJBk6WT+y3w
Q5Listnd+JEPTyDNrsj+dj3Xq3as+nCFfaWyGQMBf2cU8+gBbv78lwFl3Z6W3hs0
MYoI2t1/7w5gCPzXJPv2HaoH/xfn01jD/WkxnvaL0TOyJfx7h64tVHqlsl9QVj8X
won/DTxgW9p3HRDO13u4oG+6HzL2pCHFZRIke2gtc10cHPeBUIWpvNnxvet2LruG
odRt3ItKcvWmEyfadIZGcImTraEorrI2t8eWZsf+x4tEppPRJ660rs3YIXKuwPfQ
rf7nNq5sq1cGBZPRs4nbXGy10Z6crQKwLuMAZZ799+oTIguaBmzYBOdv4K7h1dwj
QmQGcq4Hbia7ByDBbZ2FcQbBQSGH26aU7+N770jequzf0Nc3mGCB5jyfT1CVIja6
i89eonHx+jSA3IFiurbxIWQsf38Xf5s5GM2chwsmBwCsPLuNcp4mRpTrjTHmCEJ4
7MXI/YiPWrutPxjmTD9hsbWR5nj0zAviFJHcpTknov9z0bDMAQBchOH/lF12OwxG
GJaCJ+xHYDMDj0WKdZRsSPQL6v+8DPg7G0CYLpjS5cwHP+g+JNTbWLPicWEt2dIn
Y1fWdGsTQdBVHXrpzuU1r/Pg9p52Z12MNM2O+EP/R5mC3SgmNJcM0/dls5OMbMTa
jQRd4ExIogF4x7tcqzObQhFTNVImgZk6jAUU3u/Zl88vt1qmqGnxVifMvMrplrFw
x1zVuLgkpeI63Qlxs9sXuSKnHT65ueOQzbSn7eSOBH2AS0Rlf6cHg2PYfWy9e3X4
ozSi6JpsM7Rx1VvB4LtD3Sj0ivhA6g4psxUWFJNlVNo+5l3+lM9pSl7fw7w9Djmz
l0fUIiVs2C4P44IRG4p0oah7fT+TzoNbBuK5Qxb27MyQY4lQMoHKdVO2V+kHQKv9
tbstaATkeGmCJULrX8pPxHkLKFsrdjda+uF2LMP9JIcQACSSqS4SaYCC/6kzueG/
J5IekqeonlwhdZNx+4EsQ3lrLblztlhFvUs40Zw3LmDl9bAWlUx8tx9DbQ1BqaGy
4najT694X201GvIhQB6+gEnb5Itx6JRwiZkeVdBBKUxOIE+A3bfir4jcqL/E/YKq
1QhaKm3aG+UOm6X+j5Pa3ddF6NxaMWRjnAa97qwjnSvMnUR8TLUAYbPcMCBwn86q
sVydEndLati4dcCYWlfGgMEQTycPDoXUWDUGkQj62zOJQOBdE+b5mDDZ6US9S8Kt
tdiPEE8AYCoRtFeCs0QORAZDlf6m0kDhbOjvLvxpRfSTQc1naACnyJHozls7+Bvk
ZqsngqoTOGDE+EywoeFVKJ+oR1y9GTKiJ/jXpATs2PtgopL6Rh3enO372fUctvQ3
t2ve4f4m4/XJ7QPQqICiJ7EfpN1xonQBC09IraPVRkhi8nUh7SrlaqLHd9jBOHAS
PbtLGYxIobELh3fMVnjydQxtHp2yWP2K+BXHAPblwbca3q783OvdgrlIxqdcs1aH
jPGcZZ7YboU7XcjbXEzk6PMCeCbFwjpmB8YwxeTNU6PVkCxSTyShk5xTarsdp0nT
BCAgnlNafoNZR9eVeuobwwzPLv1MPVQevIbifeHFXAJHQiEHOBV47P0VPMQkEU3o
lRWi0RhFC7VYwhe7GHZXnOlXpBSXW6wZJ650Enf8D2efR+4OV/ato55OTG1y8szN
iXuqUbmP24qn7GkZwfDf7FVI5EzD9o5Fu1FQYW7o4c2Xi/F6FeE4ZeJaCnfUZDLs
/MZjO4F/9FBuYidwAyF+LlNfTG9swSwfA0QHOT269zbhXS+UUtKAAvRNwqERNYZI
iq1sHsw1MMCV6bVSgF+YmhDWECex1eGgUaivzAEIBP1SOZmzBoO8d5JqJaGbMLB+
KXy6aW2A8gTsVOCtZdC33IaTILcRTDh+oO5LItoTTElPIfmWxVM3bLpGQU37GMOh
JYpvKmgiypnEre5H9a98v6MHBOdcmWY4+kQMiiIS+Nq16PGbKLrAP8Gw3IBa/2JA
I5J4BHRJYv/45HcHEsySKasmDbrYhNYk5GbnpydTUQmSQL3Yk9qVGhY6vTkuz4mN
B0EPh2hDyCz8qBiDhZJmclw6/c0R0FHIfn7D04KVMJe8/16P6Da7NEpieQo8m2u3
4dVl4/Mb/pX/JJL2ozVDxQezkF1N5CR1xkS4DYRbqTqoR8kQbagxLmbR1dRlDT3Q
v5YURcE69kGVcoXy9FfWRDnhdo/+3mJQr5pUxCwkUvtWvt++5xThCoACVspfiiMF
UO1o/Yb1VPvvYgXGzb7wYGD3EWxoAalAJGhmysspvAjk/+4s/nVA2WKdQoAtaSMf
DN9j/L/AN8iDxn29nEcDnevvLIcSGN4nSjuLwKkZ7NafobM6PZ8ygQIV1ACmbH06
30wlehpmrXlw9foNCNIIKtbd9uDyRNSzg+4avhyFG166Gc9OtD+sttZH2a9n+CAK
MfGdNv9mm1DNkL4Q5v0DFaULeRFRT6fxs39Nok4PBIpc6Xjw1vKo6DWXWaAxQWKi
mwlTHUCS6EBTnT59LX2CC5aYgaxlrjKOFk2VEby2HvMJLdjAQBhln7/paOPtbidb
drGCEkcdL69uNyDQBqqc8VUkILVMd4rxPimDaacP43WhzgYkPbeIqQKsAt9CPPt2
giPJ3zc/N8HNAexPWW8cweaM8wgwMsUo4Tv4nSCJl0m0leqkZZJweOI8bv1SHKct
jf9kEKojKJ013CofLcBOIJPhDAtChh6a1MFDdOq9auXOfulK2/JbCX70Rno2yvb8
mvsJTM6InukiErS2FA6wLffHLIgLTK47pTq9+mk2GLpCEFBtMZ5kZkrXKDLDc6qO
1wQFwomnFGr0aZRTXhtzVZrhTDevNOZVgREGgvnw60axmBtUZAwtwTY73wS4nxAX
flIa9miSF059A9Rz9u/vCBeb9Z0onphOquxle+C7uKhiuDl2vunq4qWpni60Pi5R
itcQnldGqjqc6tq+XgqXhmfMrvnwDv4NU2GoUF1BDM+eG1acDwqVlY4wzhpXm6I8
Y6CLtBZrLgJGS75CoU5lPbpOxn6J8hNEuKCG1SMyv54LOTLSbGPx0YGEC/H7iKs6
qmAZwYWPavuhGDdeNRYu+2AI9WEHq/7GfbEKqDWXKz0twbSZzDHBsTpkOqW6sAhY
eh6+5YDtEg8irDVH0Lp0qAZCCoR7d8w6V5VH/xl/xvZLa2RXmmVMXkA5KgGaBBKT
1vegfhYfeyKk/omefbbxKS4zSocqRS7dSB3Z0KK4qAcqgElYKoqdf/AbJx/Uk1Rg
5GcfubeO2eMaP+IZ9KTxhljc0jbozJY0buYX1skkGDzmuMhYKs6GzMtN9j78lI94
fbnrt4JN/1nCf2ea1ttJX0gf0/ab7a8GZ4fjKbkcK+aCTrZLuKkzkG5D3oc0NZ2I
1oNauuZjCqpvcN7rCLrB1C2InrRXoxjJHWeHbSKBZfwUcrAfbc4zTtpfASslKU4a
Qk80Gh4RhxfW8TYKGuVg7BFG9XMUI4WvoD/6mun534aTw6Zjq7z5URX1krSQLctr
CC9xb931H1hwDmY7l4XL/RqVROrnXJDvq23s/TDJ5lN2A3O49HhoAE6UPBe0dg5P
Wbe/P3h9cmn/m0RHKBny628SobcW6p6pM90cha7ciYSShooJ+3IzjqR6/BWFck/v
ToCK4BQ5Uicu7Is9ewY95hpMj+TyM5UtA85O2kxkQi8FMTgVdEQHpQKAuN95Gzot
sKl2HHyFUNABNNlG+ZUwCqH8WzT28wai51KiYv6ainQDMpCvsRDEUI01PgrmNkXR
8k++VX0Dj9l5aAeJ6H1vB75m31tHUsFEhiSOvbm0Vu0WW61JRIJN8wP5X3LBypKG
O5T8bPrpjLiPO+IPNzQXlvrWno8cIAwsvbvay0bIZoFCqlH+pHiU9/LIsckqgQ6m
50ub6ZadSgyP3+MegGg+RCmR56X6gI4sDDEPA7q1KGRBMr/nOmZbIMnx6MnH2/MH
zxJoCai8QURmzi5y+12vuChbahEG1NTyGOM0U8xpUpcfE0UeHCv1rNSsYft4suUV
cXHi63Pbr7tO9N5AuAuB5bRmOIc4x0bcd/+CstYN7z66F2Zmq6epGqPKcz8QfJwg
HTTwzSsozMMT8uaZDhJRBVrXGIJDkDef2e52xYzbcCkzBX3AXYfm+ziHJsnHyIUY
hY6HRjK1A+Pr8faHI2YNXg+k7tjrHVXK0DF4H3VjnhNpPVbta4xMeh7rOp4zVvOI
ur2zA3Sk7X/X9UmGUBZdJ4YoXB7nDf+GmTru8sz984ximTHjHxg1d4X0UUsqogg2
/6Ca8vtxemBG9dYZWVYZOu4M82j0cpERIHulpAgwDwgLkiOO0TsVPBafiG656/al
sHRfhH3o0fLMuYjzM9Sjp5vVSIsndaKgVavK96RW7qDA9L9lRGm8O8BXvoTp6NYi
R99NCRHxCPE0rG0VK//i5XVvGR82uPvGEyyxDMHfqv6cp2FqmyFrCZklTarmDt7l
c2o0mu5HusLu1iLCUOT5L0OKWt1TBgwAxUwLaxrJohJGMU/RpPUMc/Dg5LdvV5OH
sJKV8+mLGA+hKNo/ViOJzWoNbadLvsVo1SP+mt3GPx3PeL0E3vWrIN3ZL66129gI
YvwT/NoRJVQcekyhHlfSdomyFdM6DuMI7FQRa6/7LXpw7mu80fCsaD4BdxXIu622
R+k7yAsUFI51+VB26Z9FGRYYR8/f/4jbtrYDY+0BlAgLhXvTD9cHEZZNwHaepzOe
A2ULlB2zdBdhC3oePXC97Xh5VeAeYg+RrVz7v0E++xYOBegLayGJs1b4MuPffIeR
3hyEj7CkLj6x422C8fRexh1oLm5IwalXBWPS6ovJZ49pr4LnZQVhjYQnGhwT28HC
CNjON4ufMH9nP2TNn9+vvLWEbTVp+rtTeX43CGOxoF7CgcmB7D9waX0EvMZ9o0gL
+Xz0oqEa2RgJ7nvp6CMtUmgjHFnrHUE1kFa5rGElTQ8=
`pragma protect end_protected
